module tt_um_top_mole99 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire clknet_0_clk;
 wire net107;
 wire hsync;
 wire next_frame;
 wire next_vertical;
 wire \top_inst.background_inst.bg_select[0] ;
 wire \top_inst.background_inst.bg_select[1] ;
 wire \top_inst.background_inst.color1[0] ;
 wire \top_inst.background_inst.color1[1] ;
 wire \top_inst.background_inst.color1[2] ;
 wire \top_inst.background_inst.color1[3] ;
 wire \top_inst.background_inst.color1[4] ;
 wire \top_inst.background_inst.color1[5] ;
 wire \top_inst.background_inst.color2[0] ;
 wire \top_inst.background_inst.color2[1] ;
 wire \top_inst.background_inst.color2[2] ;
 wire \top_inst.background_inst.color2[3] ;
 wire \top_inst.background_inst.color2[4] ;
 wire \top_inst.background_inst.color2[5] ;
 wire \top_inst.background_inst.color3[0] ;
 wire \top_inst.background_inst.color3[1] ;
 wire \top_inst.background_inst.color3[2] ;
 wire \top_inst.background_inst.color3[3] ;
 wire \top_inst.background_inst.color3[4] ;
 wire \top_inst.background_inst.color3[5] ;
 wire \top_inst.background_inst.color4[0] ;
 wire \top_inst.background_inst.color4[1] ;
 wire \top_inst.background_inst.color4[2] ;
 wire \top_inst.background_inst.color4[3] ;
 wire \top_inst.background_inst.color4[4] ;
 wire \top_inst.background_inst.color4[5] ;
 wire \top_inst.background_inst.counter_h[0] ;
 wire \top_inst.background_inst.counter_h[10] ;
 wire \top_inst.background_inst.counter_h[11] ;
 wire \top_inst.background_inst.counter_h[1] ;
 wire \top_inst.background_inst.counter_h[2] ;
 wire \top_inst.background_inst.counter_h[3] ;
 wire \top_inst.background_inst.counter_h[4] ;
 wire \top_inst.background_inst.counter_h[5] ;
 wire \top_inst.background_inst.counter_h[6] ;
 wire \top_inst.background_inst.counter_h[7] ;
 wire \top_inst.background_inst.counter_h[8] ;
 wire \top_inst.background_inst.counter_h[9] ;
 wire \top_inst.background_inst.counter_v[0] ;
 wire \top_inst.background_inst.counter_v[10] ;
 wire \top_inst.background_inst.counter_v[1] ;
 wire \top_inst.background_inst.counter_v[2] ;
 wire \top_inst.background_inst.counter_v[3] ;
 wire \top_inst.background_inst.counter_v[4] ;
 wire \top_inst.background_inst.counter_v[5] ;
 wire \top_inst.background_inst.counter_v[6] ;
 wire \top_inst.background_inst.counter_v[7] ;
 wire \top_inst.background_inst.counter_v[8] ;
 wire \top_inst.background_inst.counter_v[9] ;
 wire \top_inst.background_inst.cur_time[0] ;
 wire \top_inst.background_inst.cur_time[1] ;
 wire \top_inst.background_inst.cur_time[2] ;
 wire \top_inst.background_inst.cur_time[3] ;
 wire \top_inst.background_inst.cur_time[4] ;
 wire \top_inst.background_inst.cur_time[5] ;
 wire \top_inst.background_inst.cur_time[6] ;
 wire \top_inst.background_inst.cur_time[7] ;
 wire \top_inst.misc[0] ;
 wire \top_inst.misc[1] ;
 wire \top_inst.misc[2] ;
 wire \top_inst.misc[3] ;
 wire \top_inst.spi_cs_sync ;
 wire \top_inst.spi_mosi_sync ;
 wire \top_inst.spi_receiver_inst.load_register ;
 wire \top_inst.spi_receiver_inst.reg_gclk[0] ;
 wire \top_inst.spi_receiver_inst.reg_gclk[1] ;
 wire \top_inst.spi_receiver_inst.reg_gclk[2] ;
 wire \top_inst.spi_receiver_inst.reg_gclk[3] ;
 wire \top_inst.spi_receiver_inst.reg_gclk[4] ;
 wire \top_inst.spi_receiver_inst.reg_gclk[5] ;
 wire \top_inst.spi_receiver_inst.reg_gclk[6] ;
 wire \top_inst.spi_receiver_inst.registers[4][0] ;
 wire \top_inst.spi_receiver_inst.registers[4][1] ;
 wire \top_inst.spi_receiver_inst.registers[4][2] ;
 wire \top_inst.spi_receiver_inst.registers[4][3] ;
 wire \top_inst.spi_receiver_inst.registers[4][4] ;
 wire \top_inst.spi_receiver_inst.registers[4][5] ;
 wire \top_inst.spi_receiver_inst.registers[4][6] ;
 wire \top_inst.spi_receiver_inst.registers[4][7] ;
 wire \top_inst.spi_receiver_inst.registers[5][0] ;
 wire \top_inst.spi_receiver_inst.registers[5][1] ;
 wire \top_inst.spi_receiver_inst.registers[5][2] ;
 wire \top_inst.spi_receiver_inst.registers[5][3] ;
 wire \top_inst.spi_receiver_inst.registers[5][4] ;
 wire \top_inst.spi_receiver_inst.registers[5][5] ;
 wire \top_inst.spi_receiver_inst.registers[5][6] ;
 wire \top_inst.spi_receiver_inst.registers[5][7] ;
 wire \top_inst.spi_receiver_inst.spi_cmd[0] ;
 wire \top_inst.spi_receiver_inst.spi_cmd[1] ;
 wire \top_inst.spi_receiver_inst.spi_cmd[2] ;
 wire \top_inst.spi_receiver_inst.spi_cnt[0] ;
 wire \top_inst.spi_receiver_inst.spi_cnt[1] ;
 wire \top_inst.spi_receiver_inst.spi_cnt[2] ;
 wire \top_inst.spi_receiver_inst.spi_data[0] ;
 wire \top_inst.spi_receiver_inst.spi_data[1] ;
 wire \top_inst.spi_receiver_inst.spi_data[2] ;
 wire \top_inst.spi_receiver_inst.spi_data[3] ;
 wire \top_inst.spi_receiver_inst.spi_data[4] ;
 wire \top_inst.spi_receiver_inst.spi_data[5] ;
 wire \top_inst.spi_receiver_inst.spi_data[6] ;
 wire \top_inst.spi_receiver_inst.spi_data[7] ;
 wire \top_inst.spi_receiver_inst.spi_mode ;
 wire \top_inst.spi_receiver_inst.spi_sclk ;
 wire \top_inst.spi_receiver_inst.spi_sclk_delayed ;
 wire \top_inst.sprite_access_inst.sprite_data ;
 wire \top_inst.sprite_access_inst.sprite_line[0] ;
 wire \top_inst.sprite_access_inst.sprite_line[10] ;
 wire \top_inst.sprite_access_inst.sprite_line[11] ;
 wire \top_inst.sprite_access_inst.sprite_line[1] ;
 wire \top_inst.sprite_access_inst.sprite_line[2] ;
 wire \top_inst.sprite_access_inst.sprite_line[3] ;
 wire \top_inst.sprite_access_inst.sprite_line[4] ;
 wire \top_inst.sprite_access_inst.sprite_line[5] ;
 wire \top_inst.sprite_access_inst.sprite_line[6] ;
 wire \top_inst.sprite_access_inst.sprite_line[7] ;
 wire \top_inst.sprite_access_inst.sprite_line[8] ;
 wire \top_inst.sprite_access_inst.sprite_line[9] ;
 wire \top_inst.sprite_data_inst.gclk ;
 wire \top_inst.sprite_data_inst.new_sprite_data ;
 wire \top_inst.sprite_data_inst.shiftf ;
 wire \top_inst.sprite_data_inst.sprite_data[100] ;
 wire \top_inst.sprite_data_inst.sprite_data[101] ;
 wire \top_inst.sprite_data_inst.sprite_data[102] ;
 wire \top_inst.sprite_data_inst.sprite_data[103] ;
 wire \top_inst.sprite_data_inst.sprite_data[104] ;
 wire \top_inst.sprite_data_inst.sprite_data[105] ;
 wire \top_inst.sprite_data_inst.sprite_data[106] ;
 wire \top_inst.sprite_data_inst.sprite_data[107] ;
 wire \top_inst.sprite_data_inst.sprite_data[108] ;
 wire \top_inst.sprite_data_inst.sprite_data[109] ;
 wire \top_inst.sprite_data_inst.sprite_data[10] ;
 wire \top_inst.sprite_data_inst.sprite_data[110] ;
 wire \top_inst.sprite_data_inst.sprite_data[111] ;
 wire \top_inst.sprite_data_inst.sprite_data[112] ;
 wire \top_inst.sprite_data_inst.sprite_data[113] ;
 wire \top_inst.sprite_data_inst.sprite_data[114] ;
 wire \top_inst.sprite_data_inst.sprite_data[115] ;
 wire \top_inst.sprite_data_inst.sprite_data[116] ;
 wire \top_inst.sprite_data_inst.sprite_data[117] ;
 wire \top_inst.sprite_data_inst.sprite_data[118] ;
 wire \top_inst.sprite_data_inst.sprite_data[119] ;
 wire \top_inst.sprite_data_inst.sprite_data[11] ;
 wire \top_inst.sprite_data_inst.sprite_data[120] ;
 wire \top_inst.sprite_data_inst.sprite_data[121] ;
 wire \top_inst.sprite_data_inst.sprite_data[122] ;
 wire \top_inst.sprite_data_inst.sprite_data[123] ;
 wire \top_inst.sprite_data_inst.sprite_data[124] ;
 wire \top_inst.sprite_data_inst.sprite_data[125] ;
 wire \top_inst.sprite_data_inst.sprite_data[126] ;
 wire \top_inst.sprite_data_inst.sprite_data[127] ;
 wire \top_inst.sprite_data_inst.sprite_data[128] ;
 wire \top_inst.sprite_data_inst.sprite_data[129] ;
 wire \top_inst.sprite_data_inst.sprite_data[12] ;
 wire \top_inst.sprite_data_inst.sprite_data[130] ;
 wire \top_inst.sprite_data_inst.sprite_data[131] ;
 wire \top_inst.sprite_data_inst.sprite_data[132] ;
 wire \top_inst.sprite_data_inst.sprite_data[133] ;
 wire \top_inst.sprite_data_inst.sprite_data[134] ;
 wire \top_inst.sprite_data_inst.sprite_data[135] ;
 wire \top_inst.sprite_data_inst.sprite_data[136] ;
 wire \top_inst.sprite_data_inst.sprite_data[137] ;
 wire \top_inst.sprite_data_inst.sprite_data[138] ;
 wire \top_inst.sprite_data_inst.sprite_data[139] ;
 wire \top_inst.sprite_data_inst.sprite_data[13] ;
 wire \top_inst.sprite_data_inst.sprite_data[140] ;
 wire \top_inst.sprite_data_inst.sprite_data[141] ;
 wire \top_inst.sprite_data_inst.sprite_data[142] ;
 wire \top_inst.sprite_data_inst.sprite_data[143] ;
 wire \top_inst.sprite_data_inst.sprite_data[14] ;
 wire \top_inst.sprite_data_inst.sprite_data[15] ;
 wire \top_inst.sprite_data_inst.sprite_data[16] ;
 wire \top_inst.sprite_data_inst.sprite_data[17] ;
 wire \top_inst.sprite_data_inst.sprite_data[18] ;
 wire \top_inst.sprite_data_inst.sprite_data[19] ;
 wire \top_inst.sprite_data_inst.sprite_data[1] ;
 wire \top_inst.sprite_data_inst.sprite_data[20] ;
 wire \top_inst.sprite_data_inst.sprite_data[21] ;
 wire \top_inst.sprite_data_inst.sprite_data[22] ;
 wire \top_inst.sprite_data_inst.sprite_data[23] ;
 wire \top_inst.sprite_data_inst.sprite_data[24] ;
 wire \top_inst.sprite_data_inst.sprite_data[25] ;
 wire \top_inst.sprite_data_inst.sprite_data[26] ;
 wire \top_inst.sprite_data_inst.sprite_data[27] ;
 wire \top_inst.sprite_data_inst.sprite_data[28] ;
 wire \top_inst.sprite_data_inst.sprite_data[29] ;
 wire \top_inst.sprite_data_inst.sprite_data[2] ;
 wire \top_inst.sprite_data_inst.sprite_data[30] ;
 wire \top_inst.sprite_data_inst.sprite_data[31] ;
 wire \top_inst.sprite_data_inst.sprite_data[32] ;
 wire \top_inst.sprite_data_inst.sprite_data[33] ;
 wire \top_inst.sprite_data_inst.sprite_data[34] ;
 wire \top_inst.sprite_data_inst.sprite_data[35] ;
 wire \top_inst.sprite_data_inst.sprite_data[36] ;
 wire \top_inst.sprite_data_inst.sprite_data[37] ;
 wire \top_inst.sprite_data_inst.sprite_data[38] ;
 wire \top_inst.sprite_data_inst.sprite_data[39] ;
 wire \top_inst.sprite_data_inst.sprite_data[3] ;
 wire \top_inst.sprite_data_inst.sprite_data[40] ;
 wire \top_inst.sprite_data_inst.sprite_data[41] ;
 wire \top_inst.sprite_data_inst.sprite_data[42] ;
 wire \top_inst.sprite_data_inst.sprite_data[43] ;
 wire \top_inst.sprite_data_inst.sprite_data[44] ;
 wire \top_inst.sprite_data_inst.sprite_data[45] ;
 wire \top_inst.sprite_data_inst.sprite_data[46] ;
 wire \top_inst.sprite_data_inst.sprite_data[47] ;
 wire \top_inst.sprite_data_inst.sprite_data[48] ;
 wire \top_inst.sprite_data_inst.sprite_data[49] ;
 wire \top_inst.sprite_data_inst.sprite_data[4] ;
 wire \top_inst.sprite_data_inst.sprite_data[50] ;
 wire \top_inst.sprite_data_inst.sprite_data[51] ;
 wire \top_inst.sprite_data_inst.sprite_data[52] ;
 wire \top_inst.sprite_data_inst.sprite_data[53] ;
 wire \top_inst.sprite_data_inst.sprite_data[54] ;
 wire \top_inst.sprite_data_inst.sprite_data[55] ;
 wire \top_inst.sprite_data_inst.sprite_data[56] ;
 wire \top_inst.sprite_data_inst.sprite_data[57] ;
 wire \top_inst.sprite_data_inst.sprite_data[58] ;
 wire \top_inst.sprite_data_inst.sprite_data[59] ;
 wire \top_inst.sprite_data_inst.sprite_data[5] ;
 wire \top_inst.sprite_data_inst.sprite_data[60] ;
 wire \top_inst.sprite_data_inst.sprite_data[61] ;
 wire \top_inst.sprite_data_inst.sprite_data[62] ;
 wire \top_inst.sprite_data_inst.sprite_data[63] ;
 wire \top_inst.sprite_data_inst.sprite_data[64] ;
 wire \top_inst.sprite_data_inst.sprite_data[65] ;
 wire \top_inst.sprite_data_inst.sprite_data[66] ;
 wire \top_inst.sprite_data_inst.sprite_data[67] ;
 wire \top_inst.sprite_data_inst.sprite_data[68] ;
 wire \top_inst.sprite_data_inst.sprite_data[69] ;
 wire \top_inst.sprite_data_inst.sprite_data[6] ;
 wire \top_inst.sprite_data_inst.sprite_data[70] ;
 wire \top_inst.sprite_data_inst.sprite_data[71] ;
 wire \top_inst.sprite_data_inst.sprite_data[72] ;
 wire \top_inst.sprite_data_inst.sprite_data[73] ;
 wire \top_inst.sprite_data_inst.sprite_data[74] ;
 wire \top_inst.sprite_data_inst.sprite_data[75] ;
 wire \top_inst.sprite_data_inst.sprite_data[76] ;
 wire \top_inst.sprite_data_inst.sprite_data[77] ;
 wire \top_inst.sprite_data_inst.sprite_data[78] ;
 wire \top_inst.sprite_data_inst.sprite_data[79] ;
 wire \top_inst.sprite_data_inst.sprite_data[7] ;
 wire \top_inst.sprite_data_inst.sprite_data[80] ;
 wire \top_inst.sprite_data_inst.sprite_data[81] ;
 wire \top_inst.sprite_data_inst.sprite_data[82] ;
 wire \top_inst.sprite_data_inst.sprite_data[83] ;
 wire \top_inst.sprite_data_inst.sprite_data[84] ;
 wire \top_inst.sprite_data_inst.sprite_data[85] ;
 wire \top_inst.sprite_data_inst.sprite_data[86] ;
 wire \top_inst.sprite_data_inst.sprite_data[87] ;
 wire \top_inst.sprite_data_inst.sprite_data[88] ;
 wire \top_inst.sprite_data_inst.sprite_data[89] ;
 wire \top_inst.sprite_data_inst.sprite_data[8] ;
 wire \top_inst.sprite_data_inst.sprite_data[90] ;
 wire \top_inst.sprite_data_inst.sprite_data[91] ;
 wire \top_inst.sprite_data_inst.sprite_data[92] ;
 wire \top_inst.sprite_data_inst.sprite_data[93] ;
 wire \top_inst.sprite_data_inst.sprite_data[94] ;
 wire \top_inst.sprite_data_inst.sprite_data[95] ;
 wire \top_inst.sprite_data_inst.sprite_data[96] ;
 wire \top_inst.sprite_data_inst.sprite_data[97] ;
 wire \top_inst.sprite_data_inst.sprite_data[98] ;
 wire \top_inst.sprite_data_inst.sprite_data[99] ;
 wire \top_inst.sprite_data_inst.sprite_data[9] ;
 wire \top_inst.sprite_movement_inst.divider ;
 wire \top_inst.sprite_movement_inst.sprite_x[0] ;
 wire \top_inst.sprite_movement_inst.sprite_x[1] ;
 wire \top_inst.sprite_movement_inst.sprite_x[2] ;
 wire \top_inst.sprite_movement_inst.sprite_x[3] ;
 wire \top_inst.sprite_movement_inst.sprite_x[4] ;
 wire \top_inst.sprite_movement_inst.sprite_x[5] ;
 wire \top_inst.sprite_movement_inst.sprite_x[6] ;
 wire \top_inst.sprite_movement_inst.sprite_x[7] ;
 wire \top_inst.sprite_movement_inst.sprite_x_dir ;
 wire \top_inst.sprite_movement_inst.sprite_y[0] ;
 wire \top_inst.sprite_movement_inst.sprite_y[1] ;
 wire \top_inst.sprite_movement_inst.sprite_y[2] ;
 wire \top_inst.sprite_movement_inst.sprite_y[3] ;
 wire \top_inst.sprite_movement_inst.sprite_y[4] ;
 wire \top_inst.sprite_movement_inst.sprite_y[5] ;
 wire \top_inst.sprite_movement_inst.sprite_y[6] ;
 wire \top_inst.sprite_movement_inst.sprite_y[7] ;
 wire \top_inst.sprite_movement_inst.sprite_y_dir ;
 wire \top_inst.sprite_x[0] ;
 wire \top_inst.sprite_x[1] ;
 wire \top_inst.sprite_x[2] ;
 wire \top_inst.sprite_x[3] ;
 wire \top_inst.sprite_x[4] ;
 wire \top_inst.sprite_x[5] ;
 wire \top_inst.sprite_x[6] ;
 wire \top_inst.sprite_x[7] ;
 wire \top_inst.sprite_y[0] ;
 wire \top_inst.sprite_y[1] ;
 wire \top_inst.sprite_y[2] ;
 wire \top_inst.sprite_y[3] ;
 wire \top_inst.sprite_y[4] ;
 wire \top_inst.sprite_y[5] ;
 wire \top_inst.sprite_y[6] ;
 wire \top_inst.sprite_y[7] ;
 wire \top_inst.synchronizer_spi_cs.pipe[0] ;
 wire \top_inst.synchronizer_spi_mosi.pipe[0] ;
 wire \top_inst.synchronizer_spi_sclk.pipe[0] ;
 wire \top_inst.time_dir ;
 wire \top_inst.timing_ver.sync ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_level_0_1_10_clk;
 wire clknet_level_1_1_11_clk;
 wire clknet_level_2_1_12_clk;
 wire clknet_level_3_1_13_clk;
 wire clknet_level_0_1_24_clk;
 wire clknet_level_1_1_25_clk;
 wire clknet_level_2_1_26_clk;
 wire clknet_level_3_1_27_clk;
 wire clknet_level_0_1_38_clk;
 wire clknet_level_1_1_39_clk;
 wire clknet_level_2_1_310_clk;
 wire clknet_level_3_1_311_clk;
 wire clknet_level_0_1_412_clk;
 wire clknet_level_1_1_413_clk;
 wire clknet_level_2_1_414_clk;
 wire clknet_level_3_1_415_clk;
 wire clknet_level_0_1_516_clk;
 wire clknet_level_1_1_517_clk;
 wire clknet_level_2_1_518_clk;
 wire clknet_level_3_1_519_clk;
 wire clknet_level_0_1_620_clk;
 wire clknet_level_1_1_621_clk;
 wire clknet_level_2_1_622_clk;
 wire clknet_level_3_1_623_clk;
 wire clknet_level_0_1_724_clk;
 wire clknet_level_1_1_725_clk;
 wire clknet_level_2_1_726_clk;
 wire clknet_level_3_1_727_clk;
 wire clknet_level_0_1_828_clk;
 wire clknet_level_1_1_829_clk;
 wire clknet_level_2_1_830_clk;
 wire clknet_level_3_1_831_clk;
 wire clknet_level_0_1_932_clk;
 wire clknet_level_1_1_933_clk;
 wire clknet_level_2_1_934_clk;
 wire clknet_level_3_1_935_clk;
 wire clknet_level_0_1_1036_clk;
 wire clknet_level_1_1_1037_clk;
 wire clknet_level_2_1_1038_clk;
 wire clknet_level_3_1_1039_clk;
 wire clknet_level_0_1_1140_clk;
 wire clknet_level_1_1_1141_clk;
 wire clknet_level_2_1_1142_clk;
 wire clknet_level_3_1_1143_clk;
 wire clknet_level_0_1_1244_clk;
 wire clknet_level_1_1_1245_clk;
 wire clknet_level_2_1_1246_clk;
 wire clknet_level_3_1_1247_clk;
 wire clknet_level_0_1_1348_clk;
 wire clknet_level_1_1_1349_clk;
 wire clknet_level_2_1_1350_clk;
 wire clknet_level_3_1_1351_clk;
 wire clknet_level_0_1_1452_clk;
 wire clknet_level_1_1_1453_clk;
 wire clknet_level_2_1_1454_clk;
 wire clknet_level_3_1_1455_clk;
 wire clknet_level_0_1_1556_clk;
 wire clknet_level_1_1_1557_clk;
 wire clknet_level_2_1_1558_clk;
 wire clknet_level_3_1_1559_clk;
 wire clknet_level_0_1_1660_clk;
 wire clknet_level_1_1_1661_clk;
 wire clknet_level_2_1_1662_clk;
 wire clknet_level_3_1_1663_clk;
 wire clknet_0__0021_;
 wire clknet_1_0__leaf__0021_;
 wire clknet_1_1__leaf__0021_;
 wire clknet_0__0020_;
 wire clknet_1_0__leaf__0020_;
 wire clknet_1_1__leaf__0020_;
 wire clknet_0__0019_;
 wire clknet_1_0__leaf__0019_;
 wire clknet_1_1__leaf__0019_;
 wire clknet_0__0018_;
 wire clknet_1_0__leaf__0018_;
 wire clknet_1_1__leaf__0018_;
 wire clknet_0__0017_;
 wire clknet_1_0__leaf__0017_;
 wire clknet_1_1__leaf__0017_;
 wire clknet_0__0016_;
 wire clknet_1_0__leaf__0016_;
 wire clknet_1_1__leaf__0016_;
 wire clknet_0__0015_;
 wire clknet_1_0__leaf__0015_;
 wire clknet_1_1__leaf__0015_;
 wire \clknet_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_0_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_1_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_2_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_3_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_4_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_5_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_6_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_7_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_8_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_9_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_10_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_11_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_12_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_13_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_14_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_4_15_0_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_0__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_1__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_2__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_3__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_4__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_5__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_6__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_7__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_8__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_9__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_10__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_11__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_12__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_13__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_14__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_15__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_16__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_17__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_18__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_19__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_20__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_21__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_22__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_23__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_24__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_25__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_26__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_27__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_28__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_29__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_30__leaf_top_inst.sprite_data_inst.gclk ;
 wire \clknet_5_31__leaf_top_inst.sprite_data_inst.gclk ;
 wire net167;

 sg13g2_buf_2 _1153_ (.A(\top_inst.background_inst.counter_h[11] ),
    .X(_0472_));
 sg13g2_buf_1 _1154_ (.A(\top_inst.background_inst.counter_h[9] ),
    .X(_0473_));
 sg13g2_and2_1 _1155_ (.A(_0473_),
    .B(\top_inst.background_inst.counter_h[8] ),
    .X(_0474_));
 sg13g2_buf_1 _1156_ (.A(\top_inst.background_inst.counter_h[5] ),
    .X(_0475_));
 sg13g2_buf_8 _1157_ (.A(\top_inst.background_inst.counter_h[4] ),
    .X(_0476_));
 sg13g2_inv_1 _1158_ (.Y(_0477_),
    .A(_0476_));
 sg13g2_buf_2 _1159_ (.A(\top_inst.background_inst.counter_h[2] ),
    .X(_0478_));
 sg13g2_buf_2 _1160_ (.A(\top_inst.background_inst.counter_h[1] ),
    .X(_0479_));
 sg13g2_buf_2 _1161_ (.A(\top_inst.background_inst.counter_h[0] ),
    .X(_0480_));
 sg13g2_nand4_1 _1162_ (.B(_0478_),
    .C(_0479_),
    .A(\top_inst.background_inst.counter_h[3] ),
    .Y(_0481_),
    .D(_0480_));
 sg13g2_or2_1 _1163_ (.X(_0482_),
    .B(_0481_),
    .A(_0477_));
 sg13g2_buf_2 _1164_ (.A(\top_inst.background_inst.counter_h[7] ),
    .X(_0483_));
 sg13g2_buf_1 _1165_ (.A(\top_inst.background_inst.counter_h[6] ),
    .X(_0484_));
 sg13g2_inv_1 _1166_ (.Y(_0485_),
    .A(_0038_));
 sg13g2_nor3_1 _1167_ (.A(_0483_),
    .B(net49),
    .C(_0485_),
    .Y(_0486_));
 sg13g2_o21ai_1 _1168_ (.B1(_0486_),
    .Y(_0487_),
    .A1(net50),
    .A2(_0482_));
 sg13g2_buf_1 _1169_ (.A(\top_inst.background_inst.counter_h[10] ),
    .X(_0488_));
 sg13g2_a21oi_1 _1170_ (.A1(_0474_),
    .A2(_0487_),
    .Y(_0489_),
    .B1(_0488_));
 sg13g2_or2_1 _1171_ (.X(_0490_),
    .B(_0489_),
    .A(_0472_));
 sg13g2_buf_2 _1172_ (.A(_0490_),
    .X(_0491_));
 sg13g2_inv_2 _1173_ (.Y(_0492_),
    .A(_0491_));
 sg13g2_buf_8 _1174_ (.A(\top_inst.background_inst.counter_v[5] ),
    .X(_0493_));
 sg13g2_buf_1 _1175_ (.A(_0493_),
    .X(_0494_));
 sg13g2_buf_1 _1176_ (.A(\top_inst.background_inst.counter_v[3] ),
    .X(_0495_));
 sg13g2_buf_1 _1177_ (.A(_0495_),
    .X(_0496_));
 sg13g2_buf_1 _1178_ (.A(\top_inst.background_inst.counter_v[1] ),
    .X(_0497_));
 sg13g2_buf_1 _1179_ (.A(\top_inst.background_inst.counter_v[0] ),
    .X(_0498_));
 sg13g2_buf_2 _1180_ (.A(\top_inst.background_inst.counter_v[2] ),
    .X(_0499_));
 sg13g2_and3_1 _1181_ (.X(_0500_),
    .A(net47),
    .B(_0498_),
    .C(_0499_));
 sg13g2_buf_1 _1182_ (.A(_0500_),
    .X(_0501_));
 sg13g2_buf_8 _1183_ (.A(\top_inst.background_inst.counter_v[4] ),
    .X(_0502_));
 sg13g2_o21ai_1 _1184_ (.B1(_0502_),
    .Y(_0503_),
    .A1(net35),
    .A2(_0501_));
 sg13g2_inv_1 _1185_ (.Y(_0504_),
    .A(_0503_));
 sg13g2_buf_8 _1186_ (.A(\top_inst.background_inst.counter_v[6] ),
    .X(_0505_));
 sg13g2_o21ai_1 _1187_ (.B1(net46),
    .Y(_0506_),
    .A1(net36),
    .A2(_0504_));
 sg13g2_buf_2 _1188_ (.A(\top_inst.background_inst.counter_v[7] ),
    .X(_0507_));
 sg13g2_nor2_1 _1189_ (.A(_0507_),
    .B(\top_inst.background_inst.counter_v[8] ),
    .Y(_0508_));
 sg13g2_buf_1 _1190_ (.A(\top_inst.background_inst.counter_v[9] ),
    .X(_0509_));
 sg13g2_buf_1 _1191_ (.A(\top_inst.background_inst.counter_v[10] ),
    .X(_0510_));
 sg13g2_inv_1 _1192_ (.Y(_0511_),
    .A(_0510_));
 sg13g2_nand2_1 _1193_ (.Y(_0512_),
    .A(_0509_),
    .B(_0511_));
 sg13g2_a21oi_2 _1194_ (.B1(_0512_),
    .Y(_0513_),
    .A2(_0508_),
    .A1(_0506_));
 sg13g2_and2_1 _1195_ (.A(_0492_),
    .B(_0513_),
    .X(_0514_));
 sg13g2_buf_1 _1196_ (.A(_0514_),
    .X(_0515_));
 sg13g2_buf_1 _1197_ (.A(_0515_),
    .X(next_frame));
 sg13g2_buf_1 _1198_ (.A(\top_inst.spi_receiver_inst.spi_cmd[0] ),
    .X(_0516_));
 sg13g2_buf_1 _1199_ (.A(\top_inst.spi_receiver_inst.spi_cmd[1] ),
    .X(_0517_));
 sg13g2_nand2b_1 _1200_ (.Y(_0518_),
    .B(\top_inst.spi_receiver_inst.load_register ),
    .A_N(\top_inst.spi_receiver_inst.spi_cmd[2] ));
 sg13g2_nor3_1 _1201_ (.A(_0516_),
    .B(_0517_),
    .C(_0518_),
    .Y(_0022_));
 sg13g2_nand2b_1 _1202_ (.Y(_0519_),
    .B(_0516_),
    .A_N(_0517_));
 sg13g2_nor2_1 _1203_ (.A(_0518_),
    .B(_0519_),
    .Y(_0023_));
 sg13g2_nand2b_1 _1204_ (.Y(_0520_),
    .B(_0517_),
    .A_N(_0516_));
 sg13g2_nor2_1 _1205_ (.A(_0518_),
    .B(_0520_),
    .Y(_0024_));
 sg13g2_nand2_1 _1206_ (.Y(_0521_),
    .A(_0516_),
    .B(_0517_));
 sg13g2_nor2_1 _1207_ (.A(_0518_),
    .B(_0521_),
    .Y(_0025_));
 sg13g2_nand2b_1 _1208_ (.Y(_0522_),
    .B(\top_inst.spi_receiver_inst.load_register ),
    .A_N(_0041_));
 sg13g2_nor3_1 _1209_ (.A(_0516_),
    .B(_0517_),
    .C(_0522_),
    .Y(_0026_));
 sg13g2_nor2_1 _1210_ (.A(_0519_),
    .B(_0522_),
    .Y(_0027_));
 sg13g2_nor2_1 _1211_ (.A(_0520_),
    .B(_0522_),
    .Y(_0028_));
 sg13g2_buf_1 _1212_ (.A(_0492_),
    .X(_0523_));
 sg13g2_buf_1 _1213_ (.A(net24),
    .X(next_vertical));
 sg13g2_nor2_1 _1214_ (.A(_0480_),
    .B(net23),
    .Y(_0030_));
 sg13g2_xnor2_1 _1215_ (.Y(_0524_),
    .A(_0479_),
    .B(_0480_));
 sg13g2_nor2_1 _1216_ (.A(net23),
    .B(_0524_),
    .Y(_0031_));
 sg13g2_inv_2 _1217_ (.Y(_0525_),
    .A(_0478_));
 sg13g2_nand2_1 _1218_ (.Y(_0526_),
    .A(_0479_),
    .B(_0480_));
 sg13g2_xnor2_1 _1219_ (.Y(_0527_),
    .A(_0525_),
    .B(_0526_));
 sg13g2_nor2_1 _1220_ (.A(next_vertical),
    .B(_0527_),
    .Y(_0032_));
 sg13g2_buf_1 _1221_ (.A(\top_inst.background_inst.counter_h[3] ),
    .X(_0528_));
 sg13g2_nor2_1 _1222_ (.A(_0525_),
    .B(_0526_),
    .Y(_0529_));
 sg13g2_xnor2_1 _1223_ (.Y(_0530_),
    .A(net45),
    .B(_0529_));
 sg13g2_nor2_1 _1224_ (.A(net23),
    .B(_0530_),
    .Y(_0033_));
 sg13g2_xnor2_1 _1225_ (.Y(_0531_),
    .A(_0477_),
    .B(_0481_));
 sg13g2_nor2_1 _1226_ (.A(net23),
    .B(_0531_),
    .Y(_0034_));
 sg13g2_nor2_1 _1227_ (.A(_0477_),
    .B(_0481_),
    .Y(_0532_));
 sg13g2_xnor2_1 _1228_ (.Y(_0533_),
    .A(_0485_),
    .B(_0532_));
 sg13g2_nor2_1 _1229_ (.A(next_vertical),
    .B(_0533_),
    .Y(_0035_));
 sg13g2_buf_1 _1230_ (.A(net24),
    .X(_0534_));
 sg13g2_nand2_1 _1231_ (.Y(_0535_),
    .A(net50),
    .B(_0532_));
 sg13g2_xnor2_1 _1232_ (.Y(_0536_),
    .A(_0040_),
    .B(_0535_));
 sg13g2_nor2_1 _1233_ (.A(net22),
    .B(_0536_),
    .Y(_0036_));
 sg13g2_inv_2 _1234_ (.Y(_0537_),
    .A(_0483_));
 sg13g2_nand3_1 _1235_ (.B(net49),
    .C(_0532_),
    .A(_0475_),
    .Y(_0538_));
 sg13g2_xnor2_1 _1236_ (.Y(_0539_),
    .A(_0537_),
    .B(_0538_));
 sg13g2_nor2_1 _1237_ (.A(net22),
    .B(_0539_),
    .Y(_0037_));
 sg13g2_buf_1 _1238_ (.A(net73),
    .X(_0540_));
 sg13g2_nand2b_1 _1239_ (.Y(_0011_),
    .B(net53),
    .A_N(\top_inst.spi_receiver_inst.spi_data[1] ));
 sg13g2_buf_1 _1240_ (.A(net70),
    .X(_0541_));
 sg13g2_and2_1 _1241_ (.A(_0541_),
    .B(\top_inst.spi_receiver_inst.spi_data[5] ),
    .X(_0007_));
 sg13g2_and2_1 _1242_ (.A(net52),
    .B(\top_inst.spi_receiver_inst.spi_data[6] ),
    .X(_0013_));
 sg13g2_and2_1 _1243_ (.A(net52),
    .B(\top_inst.spi_receiver_inst.spi_data[7] ),
    .X(_0014_));
 sg13g2_nand2b_1 _1244_ (.Y(_0005_),
    .B(_0540_),
    .A_N(\top_inst.spi_receiver_inst.spi_data[5] ));
 sg13g2_and2_1 _1245_ (.A(net52),
    .B(\top_inst.spi_receiver_inst.spi_data[0] ),
    .X(_0008_));
 sg13g2_nand2b_1 _1246_ (.Y(_0009_),
    .B(net53),
    .A_N(\top_inst.spi_receiver_inst.spi_data[3] ));
 sg13g2_and2_1 _1247_ (.A(_0541_),
    .B(\top_inst.spi_receiver_inst.spi_data[4] ),
    .X(_0010_));
 sg13g2_nand2b_1 _1248_ (.Y(_0006_),
    .B(net53),
    .A_N(\top_inst.spi_receiver_inst.spi_data[2] ));
 sg13g2_nand2b_1 _1249_ (.Y(_0000_),
    .B(net53),
    .A_N(\top_inst.spi_receiver_inst.spi_data[0] ));
 sg13g2_and2_1 _1250_ (.A(\top_inst.spi_receiver_inst.spi_data[1] ),
    .B(net73),
    .X(_0001_));
 sg13g2_and2_1 _1251_ (.A(net52),
    .B(\top_inst.spi_receiver_inst.spi_data[2] ),
    .X(_0002_));
 sg13g2_and2_1 _1252_ (.A(net52),
    .B(\top_inst.spi_receiver_inst.spi_data[3] ),
    .X(_0003_));
 sg13g2_nand2b_1 _1253_ (.Y(_0004_),
    .B(net53),
    .A_N(\top_inst.spi_receiver_inst.spi_data[4] ));
 sg13g2_nor2b_1 _1254_ (.A(\top_inst.spi_receiver_inst.reg_gclk[1] ),
    .B_N(_0540_),
    .Y(_0020_));
 sg13g2_nor2b_1 _1255_ (.A(\top_inst.spi_receiver_inst.reg_gclk[4] ),
    .B_N(net53),
    .Y(_0017_));
 sg13g2_inv_1 _1256_ (.Y(_0542_),
    .A(\top_inst.spi_receiver_inst.spi_cnt[2] ));
 sg13g2_inv_1 _1257_ (.Y(_0543_),
    .A(\top_inst.spi_receiver_inst.spi_sclk_delayed ));
 sg13g2_nor3_1 _1258_ (.A(_0543_),
    .B(\top_inst.spi_receiver_inst.spi_sclk ),
    .C(\top_inst.spi_cs_sync ),
    .Y(_0544_));
 sg13g2_nor2b_2 _1259_ (.A(net2),
    .B_N(_0544_),
    .Y(_0545_));
 sg13g2_nand3_1 _1260_ (.B(\top_inst.spi_receiver_inst.spi_cnt[0] ),
    .C(_0545_),
    .A(\top_inst.spi_receiver_inst.spi_cnt[1] ),
    .Y(_0546_));
 sg13g2_nor2_1 _1261_ (.A(_0542_),
    .B(_0546_),
    .Y(_0547_));
 sg13g2_and2_1 _1262_ (.A(\top_inst.spi_receiver_inst.spi_mode ),
    .B(_0547_),
    .X(_0012_));
 sg13g2_nor2b_1 _1263_ (.A(\top_inst.spi_receiver_inst.reg_gclk[3] ),
    .B_N(net53),
    .Y(_0018_));
 sg13g2_nor2b_1 _1264_ (.A(\top_inst.spi_receiver_inst.reg_gclk[6] ),
    .B_N(net53),
    .Y(_0015_));
 sg13g2_nor2b_1 _1265_ (.A(\top_inst.spi_receiver_inst.reg_gclk[2] ),
    .B_N(net52),
    .Y(_0019_));
 sg13g2_nor2b_1 _1266_ (.A(\top_inst.spi_receiver_inst.reg_gclk[0] ),
    .B_N(net52),
    .Y(_0021_));
 sg13g2_nor2b_1 _1267_ (.A(\top_inst.spi_receiver_inst.reg_gclk[5] ),
    .B_N(net52),
    .Y(_0016_));
 sg13g2_buf_1 _1268_ (.A(\top_inst.background_inst.bg_select[0] ),
    .X(_0548_));
 sg13g2_buf_1 _1269_ (.A(net44),
    .X(_0549_));
 sg13g2_nand2_1 _1270_ (.Y(_0550_),
    .A(_0523_),
    .B(_0501_));
 sg13g2_mux2_1 _1271_ (.A0(\top_inst.misc[0] ),
    .A1(net34),
    .S(_0550_),
    .X(_0102_));
 sg13g2_nand2_1 _1272_ (.Y(_0551_),
    .A(_0047_),
    .B(_0550_));
 sg13g2_o21ai_1 _1273_ (.B1(_0551_),
    .Y(_0103_),
    .A1(\top_inst.misc[1] ),
    .A2(_0550_));
 sg13g2_buf_2 _1274_ (.A(\top_inst.background_inst.cur_time[0] ),
    .X(_0552_));
 sg13g2_inv_1 _1275_ (.Y(_0553_),
    .A(_0552_));
 sg13g2_nand2_1 _1276_ (.Y(_0554_),
    .A(_0043_),
    .B(net19));
 sg13g2_o21ai_1 _1277_ (.B1(_0554_),
    .Y(_0104_),
    .A1(_0553_),
    .A2(net19));
 sg13g2_buf_1 _1278_ (.A(\top_inst.background_inst.cur_time[1] ),
    .X(_0555_));
 sg13g2_buf_2 _1279_ (.A(\top_inst.time_dir ),
    .X(_0556_));
 sg13g2_xnor2_1 _1280_ (.Y(_0557_),
    .A(_0556_),
    .B(_0043_));
 sg13g2_nand2_1 _1281_ (.Y(_0558_),
    .A(net19),
    .B(_0557_));
 sg13g2_xnor2_1 _1282_ (.Y(_0105_),
    .A(net43),
    .B(_0558_));
 sg13g2_buf_1 _1283_ (.A(\top_inst.background_inst.cur_time[2] ),
    .X(_0559_));
 sg13g2_inv_2 _1284_ (.Y(_0560_),
    .A(_0556_));
 sg13g2_a21oi_1 _1285_ (.A1(_0552_),
    .A2(_0556_),
    .Y(_0561_),
    .B1(net43));
 sg13g2_a21oi_2 _1286_ (.B1(_0561_),
    .Y(_0562_),
    .A2(_0560_),
    .A1(_0553_));
 sg13g2_xnor2_1 _1287_ (.Y(_0563_),
    .A(_0560_),
    .B(_0562_));
 sg13g2_nand2_1 _1288_ (.Y(_0564_),
    .A(net19),
    .B(_0563_));
 sg13g2_xnor2_1 _1289_ (.Y(_0106_),
    .A(net42),
    .B(_0564_));
 sg13g2_buf_1 _1290_ (.A(\top_inst.background_inst.cur_time[3] ),
    .X(_0565_));
 sg13g2_inv_2 _1291_ (.Y(_0566_),
    .A(\top_inst.background_inst.cur_time[2] ));
 sg13g2_nand2_1 _1292_ (.Y(_0567_),
    .A(_0566_),
    .B(_0556_));
 sg13g2_nand3_1 _1293_ (.B(_0560_),
    .C(_0562_),
    .A(net42),
    .Y(_0568_));
 sg13g2_o21ai_1 _1294_ (.B1(_0568_),
    .Y(_0569_),
    .A1(_0562_),
    .A2(_0567_));
 sg13g2_nand2_1 _1295_ (.Y(_0570_),
    .A(net19),
    .B(_0569_));
 sg13g2_xnor2_1 _1296_ (.Y(_0107_),
    .A(net41),
    .B(_0570_));
 sg13g2_buf_2 _1297_ (.A(\top_inst.background_inst.cur_time[4] ),
    .X(_0571_));
 sg13g2_buf_1 _1298_ (.A(_0571_),
    .X(_0572_));
 sg13g2_nand3_1 _1299_ (.B(net42),
    .C(_0562_),
    .A(net41),
    .Y(_0573_));
 sg13g2_nor2_1 _1300_ (.A(_0556_),
    .B(_0573_),
    .Y(_0574_));
 sg13g2_nor3_1 _1301_ (.A(net41),
    .B(_0562_),
    .C(_0567_),
    .Y(_0575_));
 sg13g2_o21ai_1 _1302_ (.B1(_0515_),
    .Y(_0576_),
    .A1(_0574_),
    .A2(_0575_));
 sg13g2_xnor2_1 _1303_ (.Y(_0108_),
    .A(net33),
    .B(_0576_));
 sg13g2_buf_8 _1304_ (.A(\top_inst.background_inst.cur_time[5] ),
    .X(_0577_));
 sg13g2_nand2_1 _1305_ (.Y(_0578_),
    .A(_0560_),
    .B(_0573_));
 sg13g2_or3_1 _1306_ (.A(net41),
    .B(_0559_),
    .C(_0562_),
    .X(_0579_));
 sg13g2_a22oi_1 _1307_ (.Y(_0580_),
    .B1(_0579_),
    .B2(_0556_),
    .A2(_0578_),
    .A1(net33));
 sg13g2_xnor2_1 _1308_ (.Y(_0581_),
    .A(_0556_),
    .B(_0580_));
 sg13g2_nand2_1 _1309_ (.Y(_0582_),
    .A(net19),
    .B(_0581_));
 sg13g2_xnor2_1 _1310_ (.Y(_0109_),
    .A(_0577_),
    .B(_0582_));
 sg13g2_buf_8 _1311_ (.A(\top_inst.background_inst.cur_time[6] ),
    .X(_0583_));
 sg13g2_inv_1 _1312_ (.Y(_0584_),
    .A(_0583_));
 sg13g2_nor2_1 _1313_ (.A(net40),
    .B(net33),
    .Y(_0585_));
 sg13g2_and2_1 _1314_ (.A(net40),
    .B(net33),
    .X(_0586_));
 sg13g2_a22oi_1 _1315_ (.Y(_0587_),
    .B1(_0586_),
    .B2(_0574_),
    .A2(_0585_),
    .A1(_0575_));
 sg13g2_nor2b_1 _1316_ (.A(_0587_),
    .B_N(_0515_),
    .Y(_0588_));
 sg13g2_xnor2_1 _1317_ (.Y(_0110_),
    .A(_0584_),
    .B(_0588_));
 sg13g2_inv_1 _1318_ (.Y(_0589_),
    .A(net40));
 sg13g2_nor3_1 _1319_ (.A(_0584_),
    .B(_0589_),
    .C(_0556_),
    .Y(_0590_));
 sg13g2_nor3_1 _1320_ (.A(_0583_),
    .B(_0577_),
    .C(_0560_),
    .Y(_0591_));
 sg13g2_mux2_1 _1321_ (.A0(_0590_),
    .A1(_0591_),
    .S(_0580_),
    .X(_0592_));
 sg13g2_nand2_1 _1322_ (.Y(_0593_),
    .A(_0515_),
    .B(_0592_));
 sg13g2_xnor2_1 _1323_ (.Y(_0111_),
    .A(\top_inst.background_inst.cur_time[7] ),
    .B(_0593_));
 sg13g2_nor2b_2 _1324_ (.A(\top_inst.spi_receiver_inst.spi_mode ),
    .B_N(_0545_),
    .Y(_0594_));
 sg13g2_mux2_1 _1325_ (.A0(_0516_),
    .A1(\top_inst.spi_mosi_sync ),
    .S(_0594_),
    .X(_0112_));
 sg13g2_mux2_1 _1326_ (.A0(_0517_),
    .A1(_0516_),
    .S(_0594_),
    .X(_0113_));
 sg13g2_mux2_1 _1327_ (.A0(\top_inst.spi_receiver_inst.spi_cmd[2] ),
    .A1(_0517_),
    .S(_0594_),
    .X(_0114_));
 sg13g2_mux2_1 _1328_ (.A0(\top_inst.spi_receiver_inst.spi_cnt[0] ),
    .A1(_0044_),
    .S(_0545_),
    .X(_0115_));
 sg13g2_nand2_1 _1329_ (.Y(_0595_),
    .A(\top_inst.spi_receiver_inst.spi_cnt[0] ),
    .B(_0545_));
 sg13g2_xnor2_1 _1330_ (.Y(_0116_),
    .A(\top_inst.spi_receiver_inst.spi_cnt[1] ),
    .B(_0595_));
 sg13g2_xnor2_1 _1331_ (.Y(_0117_),
    .A(\top_inst.spi_receiver_inst.spi_cnt[2] ),
    .B(_0546_));
 sg13g2_nand2_1 _1332_ (.Y(_0596_),
    .A(\top_inst.spi_receiver_inst.spi_mode ),
    .B(_0545_));
 sg13g2_buf_4 _1333_ (.X(_0597_),
    .A(_0596_));
 sg13g2_mux2_1 _1334_ (.A0(\top_inst.spi_mosi_sync ),
    .A1(\top_inst.spi_receiver_inst.spi_data[0] ),
    .S(_0597_),
    .X(_0118_));
 sg13g2_mux2_1 _1335_ (.A0(\top_inst.spi_receiver_inst.spi_data[0] ),
    .A1(\top_inst.spi_receiver_inst.spi_data[1] ),
    .S(_0597_),
    .X(_0119_));
 sg13g2_mux2_1 _1336_ (.A0(\top_inst.spi_receiver_inst.spi_data[1] ),
    .A1(\top_inst.spi_receiver_inst.spi_data[2] ),
    .S(_0597_),
    .X(_0120_));
 sg13g2_mux2_1 _1337_ (.A0(\top_inst.spi_receiver_inst.spi_data[2] ),
    .A1(\top_inst.spi_receiver_inst.spi_data[3] ),
    .S(_0597_),
    .X(_0121_));
 sg13g2_mux2_1 _1338_ (.A0(\top_inst.spi_receiver_inst.spi_data[3] ),
    .A1(\top_inst.spi_receiver_inst.spi_data[4] ),
    .S(_0597_),
    .X(_0122_));
 sg13g2_mux2_1 _1339_ (.A0(\top_inst.spi_receiver_inst.spi_data[4] ),
    .A1(\top_inst.spi_receiver_inst.spi_data[5] ),
    .S(_0597_),
    .X(_0123_));
 sg13g2_mux2_1 _1340_ (.A0(\top_inst.spi_receiver_inst.spi_data[5] ),
    .A1(\top_inst.spi_receiver_inst.spi_data[6] ),
    .S(_0597_),
    .X(_0124_));
 sg13g2_mux2_1 _1341_ (.A0(\top_inst.spi_receiver_inst.spi_data[6] ),
    .A1(\top_inst.spi_receiver_inst.spi_data[7] ),
    .S(_0597_),
    .X(_0125_));
 sg13g2_xor2_1 _1342_ (.B(_0547_),
    .A(\top_inst.spi_receiver_inst.spi_mode ),
    .X(_0126_));
 sg13g2_nand2_1 _1343_ (.Y(_0598_),
    .A(\top_inst.sprite_x[6] ),
    .B(\top_inst.sprite_x[5] ));
 sg13g2_buf_2 _1344_ (.A(\top_inst.sprite_x[3] ),
    .X(_0599_));
 sg13g2_buf_2 _1345_ (.A(\top_inst.sprite_x[2] ),
    .X(_0600_));
 sg13g2_o21ai_1 _1346_ (.B1(\top_inst.sprite_x[4] ),
    .Y(_0601_),
    .A1(_0599_),
    .A2(_0600_));
 sg13g2_buf_1 _1347_ (.A(_0601_),
    .X(_0602_));
 sg13g2_nor2_1 _1348_ (.A(_0598_),
    .B(_0602_),
    .Y(_0603_));
 sg13g2_xnor2_1 _1349_ (.Y(_0604_),
    .A(\top_inst.sprite_x[7] ),
    .B(_0603_));
 sg13g2_nand2_1 _1350_ (.Y(_0605_),
    .A(net48),
    .B(_0604_));
 sg13g2_inv_1 _1351_ (.Y(_0606_),
    .A(\top_inst.background_inst.counter_h[8] ));
 sg13g2_inv_1 _1352_ (.Y(_0607_),
    .A(\top_inst.sprite_x[5] ));
 sg13g2_nand2_1 _1353_ (.Y(_0608_),
    .A(_0607_),
    .B(_0602_));
 sg13g2_nand3_1 _1354_ (.B(\top_inst.sprite_x[6] ),
    .C(_0608_),
    .A(_0606_),
    .Y(_0609_));
 sg13g2_o21ai_1 _1355_ (.B1(\top_inst.background_inst.counter_h[8] ),
    .Y(_0610_),
    .A1(_0607_),
    .A2(_0602_));
 sg13g2_nand2_1 _1356_ (.Y(_0611_),
    .A(_0608_),
    .B(_0610_));
 sg13g2_inv_1 _1357_ (.Y(_0612_),
    .A(\top_inst.sprite_x[6] ));
 sg13g2_a221oi_1 _1358_ (.B2(_0612_),
    .C1(_0603_),
    .B1(_0611_),
    .A1(net51),
    .Y(_0613_),
    .A2(_0609_));
 sg13g2_xor2_1 _1359_ (.B(_0040_),
    .A(_0599_),
    .X(_0614_));
 sg13g2_and2_1 _1360_ (.A(net50),
    .B(_0600_),
    .X(_0615_));
 sg13g2_nand2b_1 _1361_ (.Y(_0616_),
    .B(net50),
    .A_N(_0600_));
 sg13g2_nor2_1 _1362_ (.A(_0614_),
    .B(_0616_),
    .Y(_0617_));
 sg13g2_nand2b_1 _1363_ (.Y(_0618_),
    .B(_0476_),
    .A_N(\top_inst.sprite_x[1] ));
 sg13g2_nor2b_1 _1364_ (.A(net45),
    .B_N(\top_inst.sprite_x[0] ),
    .Y(_0619_));
 sg13g2_nor2b_1 _1365_ (.A(_0476_),
    .B_N(\top_inst.sprite_x[1] ),
    .Y(_0620_));
 sg13g2_a21oi_1 _1366_ (.A1(_0618_),
    .A2(_0619_),
    .Y(_0621_),
    .B1(_0620_));
 sg13g2_a22oi_1 _1367_ (.Y(_0622_),
    .B1(_0617_),
    .B2(_0621_),
    .A2(_0615_),
    .A1(_0614_));
 sg13g2_and2_1 _1368_ (.A(_0600_),
    .B(_0614_),
    .X(_0623_));
 sg13g2_or3_1 _1369_ (.A(_0599_),
    .B(_0600_),
    .C(\top_inst.sprite_x[4] ),
    .X(_0624_));
 sg13g2_nand2_1 _1370_ (.Y(_0625_),
    .A(_0602_),
    .B(_0624_));
 sg13g2_xor2_1 _1371_ (.B(_0600_),
    .A(_0599_),
    .X(_0626_));
 sg13g2_and2_1 _1372_ (.A(net49),
    .B(_0626_),
    .X(_0627_));
 sg13g2_a221oi_1 _1373_ (.B2(_0483_),
    .C1(_0627_),
    .B1(_0625_),
    .A1(_0623_),
    .Y(_0628_),
    .A2(_0621_));
 sg13g2_nor2_1 _1374_ (.A(_0483_),
    .B(_0625_),
    .Y(_0629_));
 sg13g2_a21o_1 _1375_ (.A2(_0628_),
    .A1(_0622_),
    .B1(_0629_),
    .X(_0630_));
 sg13g2_or2_1 _1376_ (.X(_0631_),
    .B(_0602_),
    .A(_0607_));
 sg13g2_xnor2_1 _1377_ (.Y(_0632_),
    .A(_0612_),
    .B(_0631_));
 sg13g2_a21oi_1 _1378_ (.A1(_0631_),
    .A2(_0608_),
    .Y(_0633_),
    .B1(_0606_));
 sg13g2_a221oi_1 _1379_ (.B2(net51),
    .C1(_0633_),
    .B1(_0632_),
    .A1(net48),
    .Y(_0634_),
    .A2(_0604_));
 sg13g2_inv_1 _1380_ (.Y(_0635_),
    .A(\top_inst.sprite_x[7] ));
 sg13g2_or3_1 _1381_ (.A(_0635_),
    .B(_0598_),
    .C(_0602_),
    .X(_0636_));
 sg13g2_or2_1 _1382_ (.X(_0637_),
    .B(_0636_),
    .A(_0472_));
 sg13g2_o21ai_1 _1383_ (.B1(_0637_),
    .Y(_0638_),
    .A1(net48),
    .A2(_0604_));
 sg13g2_a221oi_1 _1384_ (.B2(_0634_),
    .C1(_0638_),
    .B1(_0630_),
    .A1(_0605_),
    .Y(_0639_),
    .A2(_0613_));
 sg13g2_inv_1 _1385_ (.Y(_0640_),
    .A(_0509_));
 sg13g2_inv_1 _1386_ (.Y(_0641_),
    .A(\top_inst.sprite_y[6] ));
 sg13g2_buf_1 _1387_ (.A(\top_inst.sprite_y[5] ),
    .X(_0642_));
 sg13g2_inv_1 _1388_ (.Y(_0643_),
    .A(_0642_));
 sg13g2_buf_1 _1389_ (.A(\top_inst.sprite_y[3] ),
    .X(_0644_));
 sg13g2_buf_2 _1390_ (.A(\top_inst.sprite_y[2] ),
    .X(_0645_));
 sg13g2_buf_2 _1391_ (.A(\top_inst.sprite_y[4] ),
    .X(_0646_));
 sg13g2_o21ai_1 _1392_ (.B1(_0646_),
    .Y(_0647_),
    .A1(_0644_),
    .A2(_0645_));
 sg13g2_nor2_1 _1393_ (.A(_0643_),
    .B(_0647_),
    .Y(_0648_));
 sg13g2_xnor2_1 _1394_ (.Y(_0649_),
    .A(_0641_),
    .B(_0648_));
 sg13g2_nand2b_1 _1395_ (.Y(_0650_),
    .B(\top_inst.sprite_y[1] ),
    .A_N(_0502_));
 sg13g2_nand2b_1 _1396_ (.Y(_0651_),
    .B(\top_inst.sprite_y[0] ),
    .A_N(net35));
 sg13g2_nor2b_1 _1397_ (.A(\top_inst.sprite_y[1] ),
    .B_N(_0502_),
    .Y(_0652_));
 sg13g2_a21oi_1 _1398_ (.A1(_0650_),
    .A2(_0651_),
    .Y(_0653_),
    .B1(_0652_));
 sg13g2_nand2_1 _1399_ (.Y(_0654_),
    .A(net36),
    .B(_0645_));
 sg13g2_xor2_1 _1400_ (.B(_0645_),
    .A(_0644_),
    .X(_0655_));
 sg13g2_or2_1 _1401_ (.X(_0656_),
    .B(_0645_),
    .A(_0493_));
 sg13g2_o21ai_1 _1402_ (.B1(_0656_),
    .Y(_0657_),
    .A1(net46),
    .A2(_0655_));
 sg13g2_a21o_1 _1403_ (.A2(_0654_),
    .A1(_0653_),
    .B1(_0657_),
    .X(_0658_));
 sg13g2_xnor2_1 _1404_ (.Y(_0659_),
    .A(_0643_),
    .B(_0647_));
 sg13g2_buf_1 _1405_ (.A(\top_inst.background_inst.counter_v[8] ),
    .X(_0660_));
 sg13g2_or3_1 _1406_ (.A(_0644_),
    .B(_0645_),
    .C(_0646_),
    .X(_0661_));
 sg13g2_inv_1 _1407_ (.Y(_0662_),
    .A(_0507_));
 sg13g2_a21oi_1 _1408_ (.A1(_0647_),
    .A2(_0661_),
    .Y(_0663_),
    .B1(_0662_));
 sg13g2_a221oi_1 _1409_ (.B2(net39),
    .C1(_0663_),
    .B1(_0659_),
    .A1(net46),
    .Y(_0664_),
    .A2(_0655_));
 sg13g2_nor2b_1 _1410_ (.A(net39),
    .B_N(_0646_),
    .Y(_0665_));
 sg13g2_or2_1 _1411_ (.X(_0666_),
    .B(_0645_),
    .A(_0644_));
 sg13g2_o21ai_1 _1412_ (.B1(_0666_),
    .Y(_0667_),
    .A1(_0508_),
    .A2(_0665_));
 sg13g2_a21oi_1 _1413_ (.A1(_0646_),
    .A2(_0508_),
    .Y(_0668_),
    .B1(_0642_));
 sg13g2_nand2_1 _1414_ (.Y(_0669_),
    .A(_0662_),
    .B(_0661_));
 sg13g2_a221oi_1 _1415_ (.B2(net39),
    .C1(_0648_),
    .B1(_0669_),
    .A1(_0667_),
    .Y(_0670_),
    .A2(_0668_));
 sg13g2_a221oi_1 _1416_ (.B2(_0664_),
    .C1(_0670_),
    .B1(_0658_),
    .A1(_0640_),
    .Y(_0671_),
    .A2(_0649_));
 sg13g2_inv_1 _1417_ (.Y(_0672_),
    .A(\top_inst.sprite_y[7] ));
 sg13g2_nand2_1 _1418_ (.Y(_0673_),
    .A(_0510_),
    .B(_0672_));
 sg13g2_o21ai_1 _1419_ (.B1(_0641_),
    .Y(_0674_),
    .A1(_0643_),
    .A2(_0647_));
 sg13g2_nor2_1 _1420_ (.A(_0511_),
    .B(\top_inst.sprite_y[7] ),
    .Y(_0675_));
 sg13g2_nand4_1 _1421_ (.B(_0642_),
    .C(_0646_),
    .A(\top_inst.sprite_y[6] ),
    .Y(_0676_),
    .D(_0666_));
 sg13g2_nand2_1 _1422_ (.Y(_0677_),
    .A(_0675_),
    .B(_0676_));
 sg13g2_a22oi_1 _1423_ (.Y(_0678_),
    .B1(_0677_),
    .B2(_0640_),
    .A2(_0674_),
    .A1(_0673_));
 sg13g2_a21oi_1 _1424_ (.A1(_0672_),
    .A2(_0676_),
    .Y(_0679_),
    .B1(_0510_));
 sg13g2_or2_1 _1425_ (.X(_0680_),
    .B(_0676_),
    .A(_0672_));
 sg13g2_nor2b_1 _1426_ (.A(_0679_),
    .B_N(_0680_),
    .Y(_0681_));
 sg13g2_o21ai_1 _1427_ (.B1(_0681_),
    .Y(_0682_),
    .A1(_0671_),
    .A2(_0678_));
 sg13g2_nand2b_1 _1428_ (.Y(_0683_),
    .B(\top_inst.sprite_x[7] ),
    .A_N(net48));
 sg13g2_nand2b_1 _1429_ (.Y(_0684_),
    .B(net49),
    .A_N(_0599_));
 sg13g2_nand3b_1 _1430_ (.B(_0683_),
    .C(_0684_),
    .Y(_0685_),
    .A_N(_0619_));
 sg13g2_nand2b_1 _1431_ (.Y(_0686_),
    .B(net45),
    .A_N(\top_inst.sprite_x[0] ));
 sg13g2_nand2b_1 _1432_ (.Y(_0687_),
    .B(\top_inst.sprite_x[6] ),
    .A_N(net51));
 sg13g2_nand4_1 _1433_ (.B(_0616_),
    .C(_0686_),
    .A(_0618_),
    .Y(_0688_),
    .D(_0687_));
 sg13g2_nand2b_1 _1434_ (.Y(_0689_),
    .B(_0483_),
    .A_N(\top_inst.sprite_x[4] ));
 sg13g2_nand2b_1 _1435_ (.Y(_0690_),
    .B(net51),
    .A_N(\top_inst.sprite_x[6] ));
 sg13g2_nand2b_1 _1436_ (.Y(_0691_),
    .B(\top_inst.sprite_x[5] ),
    .A_N(\top_inst.background_inst.counter_h[8] ));
 sg13g2_nand2b_1 _1437_ (.Y(_0692_),
    .B(\top_inst.background_inst.counter_h[8] ),
    .A_N(\top_inst.sprite_x[5] ));
 sg13g2_nand4_1 _1438_ (.B(_0690_),
    .C(_0691_),
    .A(_0689_),
    .Y(_0693_),
    .D(_0692_));
 sg13g2_nor2b_1 _1439_ (.A(_0483_),
    .B_N(\top_inst.sprite_x[4] ),
    .Y(_0694_));
 sg13g2_nor2b_1 _1440_ (.A(net49),
    .B_N(_0599_),
    .Y(_0695_));
 sg13g2_nor2b_1 _1441_ (.A(net50),
    .B_N(_0600_),
    .Y(_0696_));
 sg13g2_or4_1 _1442_ (.A(_0620_),
    .B(_0694_),
    .C(_0695_),
    .D(_0696_),
    .X(_0697_));
 sg13g2_nor4_1 _1443_ (.A(_0685_),
    .B(_0688_),
    .C(_0693_),
    .D(_0697_),
    .Y(_0698_));
 sg13g2_a21oi_1 _1444_ (.A1(net48),
    .A2(_0635_),
    .Y(_0699_),
    .B1(_0472_));
 sg13g2_nor2b_1 _1445_ (.A(_0698_),
    .B_N(_0699_),
    .Y(_0700_));
 sg13g2_nand2_1 _1446_ (.Y(_0701_),
    .A(_0618_),
    .B(_0686_));
 sg13g2_nor4_1 _1447_ (.A(_0620_),
    .B(_0694_),
    .C(_0695_),
    .D(_0696_),
    .Y(_0702_));
 sg13g2_o21ai_1 _1448_ (.B1(_0684_),
    .Y(_0703_),
    .A1(_0616_),
    .A2(_0695_));
 sg13g2_nand2_1 _1449_ (.Y(_0704_),
    .A(_0537_),
    .B(\top_inst.sprite_x[4] ));
 sg13g2_a221oi_1 _1450_ (.B2(_0704_),
    .C1(_0693_),
    .B1(_0703_),
    .A1(_0701_),
    .Y(_0705_),
    .A2(_0702_));
 sg13g2_inv_1 _1451_ (.Y(_0706_),
    .A(net48));
 sg13g2_o21ai_1 _1452_ (.B1(_0612_),
    .Y(_0707_),
    .A1(net51),
    .A2(_0691_));
 sg13g2_nand2_1 _1453_ (.Y(_0708_),
    .A(net51),
    .B(_0691_));
 sg13g2_a22oi_1 _1454_ (.Y(_0709_),
    .B1(_0707_),
    .B2(_0708_),
    .A2(\top_inst.sprite_x[7] ),
    .A1(_0706_));
 sg13g2_nand2b_1 _1455_ (.Y(_0710_),
    .B(_0709_),
    .A_N(_0705_));
 sg13g2_nand2_1 _1456_ (.Y(_0711_),
    .A(net39),
    .B(_0643_));
 sg13g2_nand2_1 _1457_ (.Y(_0712_),
    .A(_0509_),
    .B(_0641_));
 sg13g2_nand4_1 _1458_ (.B(_0646_),
    .C(_0711_),
    .A(_0662_),
    .Y(_0713_),
    .D(_0712_));
 sg13g2_nand2_1 _1459_ (.Y(_0714_),
    .A(_0640_),
    .B(\top_inst.sprite_y[6] ));
 sg13g2_nand3b_1 _1460_ (.B(_0642_),
    .C(_0712_),
    .Y(_0715_),
    .A_N(net39));
 sg13g2_nand3_1 _1461_ (.B(_0714_),
    .C(_0715_),
    .A(_0713_),
    .Y(_0716_));
 sg13g2_inv_1 _1462_ (.Y(_0717_),
    .A(_0644_));
 sg13g2_xor2_1 _1463_ (.B(_0642_),
    .A(net39),
    .X(_0718_));
 sg13g2_a221oi_1 _1464_ (.B2(_0510_),
    .C1(_0718_),
    .B1(_0672_),
    .A1(net46),
    .Y(_0719_),
    .A2(_0717_));
 sg13g2_xnor2_1 _1465_ (.Y(_0720_),
    .A(_0507_),
    .B(_0646_));
 sg13g2_nand4_1 _1466_ (.B(_0714_),
    .C(_0719_),
    .A(_0712_),
    .Y(_0721_),
    .D(_0720_));
 sg13g2_inv_1 _1467_ (.Y(_0722_),
    .A(_0505_));
 sg13g2_inv_1 _1468_ (.Y(_0723_),
    .A(_0645_));
 sg13g2_nand2_1 _1469_ (.Y(_0724_),
    .A(net36),
    .B(_0723_));
 sg13g2_nor2_1 _1470_ (.A(net36),
    .B(_0723_),
    .Y(_0725_));
 sg13g2_a221oi_1 _1471_ (.B2(_0653_),
    .C1(_0725_),
    .B1(_0724_),
    .A1(_0722_),
    .Y(_0726_),
    .A2(_0644_));
 sg13g2_a22oi_1 _1472_ (.Y(_0727_),
    .B1(_0636_),
    .B2(_0472_),
    .A2(\top_inst.sprite_y[7] ),
    .A1(_0511_));
 sg13g2_o21ai_1 _1473_ (.B1(_0727_),
    .Y(_0728_),
    .A1(_0721_),
    .A2(_0726_));
 sg13g2_a221oi_1 _1474_ (.B2(_0716_),
    .C1(_0728_),
    .B1(_0673_),
    .A1(_0700_),
    .Y(_0729_),
    .A2(_0710_));
 sg13g2_nand3b_1 _1475_ (.B(_0682_),
    .C(_0729_),
    .Y(_0730_),
    .A_N(_0639_));
 sg13g2_buf_2 _1476_ (.A(_0730_),
    .X(_0731_));
 sg13g2_nor3_2 _1477_ (.A(_0525_),
    .B(_0526_),
    .C(_0731_),
    .Y(_0732_));
 sg13g2_buf_1 _1478_ (.A(_0732_),
    .X(_0733_));
 sg13g2_buf_1 _1479_ (.A(_0498_),
    .X(_0734_));
 sg13g2_buf_1 _1480_ (.A(_0499_),
    .X(_0735_));
 sg13g2_nor3_1 _1481_ (.A(net47),
    .B(_0734_),
    .C(_0735_),
    .Y(_0736_));
 sg13g2_mux2_1 _1482_ (.A0(\top_inst.sprite_access_inst.sprite_line[11] ),
    .A1(\top_inst.sprite_access_inst.sprite_data ),
    .S(_0736_),
    .X(_0737_));
 sg13g2_inv_1 _1483_ (.Y(_0738_),
    .A(_0737_));
 sg13g2_buf_1 _1484_ (.A(_0738_),
    .X(_0739_));
 sg13g2_nor2_1 _1485_ (.A(\top_inst.sprite_access_inst.sprite_line[0] ),
    .B(net18),
    .Y(_0740_));
 sg13g2_a21oi_1 _1486_ (.A1(net18),
    .A2(_0739_),
    .Y(_0127_),
    .B1(_0740_));
 sg13g2_mux2_1 _1487_ (.A0(\top_inst.sprite_access_inst.sprite_line[10] ),
    .A1(\top_inst.sprite_access_inst.sprite_line[9] ),
    .S(net18),
    .X(_0128_));
 sg13g2_mux2_1 _1488_ (.A0(\top_inst.sprite_access_inst.sprite_line[11] ),
    .A1(\top_inst.sprite_access_inst.sprite_line[10] ),
    .S(net18),
    .X(_0129_));
 sg13g2_mux2_1 _1489_ (.A0(\top_inst.sprite_access_inst.sprite_line[1] ),
    .A1(\top_inst.sprite_access_inst.sprite_line[0] ),
    .S(net18),
    .X(_0130_));
 sg13g2_mux2_1 _1490_ (.A0(\top_inst.sprite_access_inst.sprite_line[2] ),
    .A1(\top_inst.sprite_access_inst.sprite_line[1] ),
    .S(_0733_),
    .X(_0131_));
 sg13g2_mux2_1 _1491_ (.A0(\top_inst.sprite_access_inst.sprite_line[3] ),
    .A1(\top_inst.sprite_access_inst.sprite_line[2] ),
    .S(_0733_),
    .X(_0132_));
 sg13g2_mux2_1 _1492_ (.A0(\top_inst.sprite_access_inst.sprite_line[4] ),
    .A1(\top_inst.sprite_access_inst.sprite_line[3] ),
    .S(net18),
    .X(_0133_));
 sg13g2_mux2_1 _1493_ (.A0(\top_inst.sprite_access_inst.sprite_line[5] ),
    .A1(\top_inst.sprite_access_inst.sprite_line[4] ),
    .S(net18),
    .X(_0134_));
 sg13g2_mux2_1 _1494_ (.A0(\top_inst.sprite_access_inst.sprite_line[6] ),
    .A1(\top_inst.sprite_access_inst.sprite_line[5] ),
    .S(_0732_),
    .X(_0135_));
 sg13g2_mux2_1 _1495_ (.A0(\top_inst.sprite_access_inst.sprite_line[7] ),
    .A1(\top_inst.sprite_access_inst.sprite_line[6] ),
    .S(_0732_),
    .X(_0136_));
 sg13g2_mux2_1 _1496_ (.A0(\top_inst.sprite_access_inst.sprite_line[8] ),
    .A1(\top_inst.sprite_access_inst.sprite_line[7] ),
    .S(_0732_),
    .X(_0137_));
 sg13g2_mux2_1 _1497_ (.A0(\top_inst.sprite_access_inst.sprite_line[9] ),
    .A1(\top_inst.sprite_access_inst.sprite_line[8] ),
    .S(_0732_),
    .X(_0138_));
 sg13g2_mux2_1 _1498_ (.A0(\top_inst.sprite_movement_inst.divider ),
    .A1(_0029_),
    .S(net19),
    .X(_0139_));
 sg13g2_buf_2 _1499_ (.A(\top_inst.sprite_movement_inst.sprite_x[0] ),
    .X(_0741_));
 sg13g2_nand3_1 _1500_ (.B(\top_inst.sprite_movement_inst.divider ),
    .C(_0515_),
    .A(\top_inst.misc[2] ),
    .Y(_0742_));
 sg13g2_buf_1 _1501_ (.A(_0742_),
    .X(_0743_));
 sg13g2_buf_1 _1502_ (.A(net17),
    .X(_0744_));
 sg13g2_mux2_1 _1503_ (.A0(_0045_),
    .A1(_0741_),
    .S(net16),
    .X(_0140_));
 sg13g2_buf_1 _1504_ (.A(\top_inst.sprite_movement_inst.sprite_x[1] ),
    .X(_0745_));
 sg13g2_inv_1 _1505_ (.Y(_0746_),
    .A(_0745_));
 sg13g2_buf_2 _1506_ (.A(\top_inst.sprite_movement_inst.sprite_x_dir ),
    .X(_0747_));
 sg13g2_xor2_1 _1507_ (.B(_0045_),
    .A(_0747_),
    .X(_0748_));
 sg13g2_nor2_1 _1508_ (.A(net16),
    .B(_0748_),
    .Y(_0749_));
 sg13g2_xnor2_1 _1509_ (.Y(_0141_),
    .A(_0746_),
    .B(_0749_));
 sg13g2_buf_2 _1510_ (.A(\top_inst.sprite_movement_inst.sprite_x[2] ),
    .X(_0750_));
 sg13g2_nor2b_1 _1511_ (.A(_0747_),
    .B_N(_0741_),
    .Y(_0751_));
 sg13g2_inv_1 _1512_ (.Y(_0752_),
    .A(_0747_));
 sg13g2_nor3_1 _1513_ (.A(_0745_),
    .B(_0741_),
    .C(_0752_),
    .Y(_0753_));
 sg13g2_a21oi_1 _1514_ (.A1(_0745_),
    .A2(_0751_),
    .Y(_0754_),
    .B1(_0753_));
 sg13g2_nor2_1 _1515_ (.A(net16),
    .B(_0754_),
    .Y(_0755_));
 sg13g2_xor2_1 _1516_ (.B(_0755_),
    .A(_0750_),
    .X(_0142_));
 sg13g2_buf_1 _1517_ (.A(\top_inst.sprite_movement_inst.sprite_x[3] ),
    .X(_0756_));
 sg13g2_and3_1 _1518_ (.X(_0757_),
    .A(_0745_),
    .B(_0750_),
    .C(_0751_));
 sg13g2_nor3_1 _1519_ (.A(_0745_),
    .B(_0741_),
    .C(_0750_),
    .Y(_0758_));
 sg13g2_nand2_1 _1520_ (.Y(_0759_),
    .A(_0747_),
    .B(_0758_));
 sg13g2_nor2b_1 _1521_ (.A(_0757_),
    .B_N(_0759_),
    .Y(_0760_));
 sg13g2_nor2_1 _1522_ (.A(_0744_),
    .B(_0760_),
    .Y(_0761_));
 sg13g2_xor2_1 _1523_ (.B(_0761_),
    .A(net38),
    .X(_0143_));
 sg13g2_buf_1 _1524_ (.A(\top_inst.sprite_movement_inst.sprite_x[4] ),
    .X(_0762_));
 sg13g2_nor2_1 _1525_ (.A(net38),
    .B(_0759_),
    .Y(_0763_));
 sg13g2_a21oi_1 _1526_ (.A1(net38),
    .A2(_0757_),
    .Y(_0764_),
    .B1(_0763_));
 sg13g2_nor2_1 _1527_ (.A(_0744_),
    .B(_0764_),
    .Y(_0765_));
 sg13g2_xor2_1 _1528_ (.B(_0765_),
    .A(net37),
    .X(_0144_));
 sg13g2_buf_2 _1529_ (.A(\top_inst.sprite_movement_inst.sprite_x[5] ),
    .X(_0766_));
 sg13g2_nand4_1 _1530_ (.B(net38),
    .C(_0750_),
    .A(_0741_),
    .Y(_0767_),
    .D(net37));
 sg13g2_or4_1 _1531_ (.A(_0741_),
    .B(net38),
    .C(_0750_),
    .D(net37),
    .X(_0768_));
 sg13g2_a21oi_1 _1532_ (.A1(_0747_),
    .A2(_0768_),
    .Y(_0769_),
    .B1(_0745_));
 sg13g2_a21oi_1 _1533_ (.A1(_0752_),
    .A2(_0767_),
    .Y(_0770_),
    .B1(_0769_));
 sg13g2_xnor2_1 _1534_ (.Y(_0771_),
    .A(_0747_),
    .B(_0770_));
 sg13g2_nor2_1 _1535_ (.A(net16),
    .B(_0771_),
    .Y(_0772_));
 sg13g2_xor2_1 _1536_ (.B(_0772_),
    .A(_0766_),
    .X(_0145_));
 sg13g2_buf_1 _1537_ (.A(\top_inst.sprite_movement_inst.sprite_x[6] ),
    .X(_0773_));
 sg13g2_or4_1 _1538_ (.A(net38),
    .B(_0766_),
    .C(net37),
    .D(_0759_),
    .X(_0774_));
 sg13g2_nand4_1 _1539_ (.B(_0766_),
    .C(net37),
    .A(net38),
    .Y(_0775_),
    .D(_0757_));
 sg13g2_a21oi_1 _1540_ (.A1(_0774_),
    .A2(_0775_),
    .Y(_0776_),
    .B1(net17));
 sg13g2_xor2_1 _1541_ (.B(_0776_),
    .A(_0773_),
    .X(_0146_));
 sg13g2_nand4_1 _1542_ (.B(_0773_),
    .C(_0752_),
    .A(_0766_),
    .Y(_0777_),
    .D(_0770_));
 sg13g2_or4_1 _1543_ (.A(_0766_),
    .B(_0773_),
    .C(_0752_),
    .D(_0770_),
    .X(_0778_));
 sg13g2_a21oi_1 _1544_ (.A1(_0777_),
    .A2(_0778_),
    .Y(_0779_),
    .B1(net17));
 sg13g2_xor2_1 _1545_ (.B(_0779_),
    .A(\top_inst.sprite_movement_inst.sprite_x[7] ),
    .X(_0147_));
 sg13g2_nand2b_1 _1546_ (.Y(_0780_),
    .B(_0741_),
    .A_N(\top_inst.sprite_movement_inst.sprite_x[7] ));
 sg13g2_nor4_1 _1547_ (.A(net38),
    .B(_0766_),
    .C(net17),
    .D(_0780_),
    .Y(_0781_));
 sg13g2_and3_1 _1548_ (.X(_0782_),
    .A(_0750_),
    .B(net37),
    .C(_0773_));
 sg13g2_a21oi_1 _1549_ (.A1(_0781_),
    .A2(_0782_),
    .Y(_0783_),
    .B1(_0747_));
 sg13g2_nor3_1 _1550_ (.A(_0750_),
    .B(net37),
    .C(_0773_),
    .Y(_0784_));
 sg13g2_a21o_1 _1551_ (.A2(_0784_),
    .A1(_0781_),
    .B1(_0752_),
    .X(_0785_));
 sg13g2_o21ai_1 _1552_ (.B1(_0785_),
    .Y(_0148_),
    .A1(_0746_),
    .A2(_0783_));
 sg13g2_buf_2 _1553_ (.A(\top_inst.sprite_movement_inst.sprite_y[0] ),
    .X(_0786_));
 sg13g2_mux2_1 _1554_ (.A0(_0046_),
    .A1(_0786_),
    .S(net16),
    .X(_0149_));
 sg13g2_buf_2 _1555_ (.A(\top_inst.sprite_movement_inst.sprite_y[1] ),
    .X(_0787_));
 sg13g2_buf_2 _1556_ (.A(\top_inst.sprite_movement_inst.sprite_y_dir ),
    .X(_0788_));
 sg13g2_xor2_1 _1557_ (.B(_0046_),
    .A(_0788_),
    .X(_0789_));
 sg13g2_nor2_1 _1558_ (.A(net16),
    .B(_0789_),
    .Y(_0790_));
 sg13g2_xor2_1 _1559_ (.B(_0790_),
    .A(_0787_),
    .X(_0150_));
 sg13g2_buf_1 _1560_ (.A(\top_inst.sprite_movement_inst.sprite_y[2] ),
    .X(_0791_));
 sg13g2_inv_1 _1561_ (.Y(_0792_),
    .A(_0791_));
 sg13g2_inv_2 _1562_ (.Y(_0793_),
    .A(_0788_));
 sg13g2_and2_1 _1563_ (.A(_0787_),
    .B(_0786_),
    .X(_0794_));
 sg13g2_nor3_2 _1564_ (.A(_0787_),
    .B(_0786_),
    .C(_0793_),
    .Y(_0795_));
 sg13g2_a21oi_1 _1565_ (.A1(_0793_),
    .A2(_0794_),
    .Y(_0796_),
    .B1(_0795_));
 sg13g2_nor2_1 _1566_ (.A(net16),
    .B(_0796_),
    .Y(_0797_));
 sg13g2_xnor2_1 _1567_ (.Y(_0151_),
    .A(_0792_),
    .B(_0797_));
 sg13g2_buf_2 _1568_ (.A(\top_inst.sprite_movement_inst.sprite_y[3] ),
    .X(_0798_));
 sg13g2_and3_1 _1569_ (.X(_0799_),
    .A(_0791_),
    .B(_0793_),
    .C(_0794_));
 sg13g2_a21oi_1 _1570_ (.A1(_0792_),
    .A2(_0795_),
    .Y(_0800_),
    .B1(_0799_));
 sg13g2_nor2_1 _1571_ (.A(net17),
    .B(_0800_),
    .Y(_0801_));
 sg13g2_xor2_1 _1572_ (.B(_0801_),
    .A(_0798_),
    .X(_0152_));
 sg13g2_buf_1 _1573_ (.A(\top_inst.sprite_movement_inst.sprite_y[4] ),
    .X(_0802_));
 sg13g2_nor2_1 _1574_ (.A(_0798_),
    .B(_0791_),
    .Y(_0803_));
 sg13g2_a22oi_1 _1575_ (.Y(_0804_),
    .B1(_0803_),
    .B2(_0795_),
    .A2(_0799_),
    .A1(_0798_));
 sg13g2_nor2_1 _1576_ (.A(net17),
    .B(_0804_),
    .Y(_0805_));
 sg13g2_xor2_1 _1577_ (.B(_0805_),
    .A(_0802_),
    .X(_0153_));
 sg13g2_buf_2 _1578_ (.A(\top_inst.sprite_movement_inst.sprite_y[5] ),
    .X(_0806_));
 sg13g2_nor4_1 _1579_ (.A(_0786_),
    .B(_0798_),
    .C(_0791_),
    .D(_0802_),
    .Y(_0807_));
 sg13g2_and4_1 _1580_ (.A(_0786_),
    .B(_0798_),
    .C(_0791_),
    .D(_0802_),
    .X(_0808_));
 sg13g2_o21ai_1 _1581_ (.B1(_0787_),
    .Y(_0809_),
    .A1(_0788_),
    .A2(_0808_));
 sg13g2_o21ai_1 _1582_ (.B1(_0809_),
    .Y(_0810_),
    .A1(_0793_),
    .A2(_0807_));
 sg13g2_xnor2_1 _1583_ (.Y(_0811_),
    .A(_0788_),
    .B(_0810_));
 sg13g2_nor2_1 _1584_ (.A(net17),
    .B(_0811_),
    .Y(_0812_));
 sg13g2_xor2_1 _1585_ (.B(_0812_),
    .A(_0806_),
    .X(_0154_));
 sg13g2_nor4_1 _1586_ (.A(_0798_),
    .B(_0791_),
    .C(_0802_),
    .D(_0806_),
    .Y(_0813_));
 sg13g2_nand2_1 _1587_ (.Y(_0814_),
    .A(_0795_),
    .B(_0813_));
 sg13g2_nand4_1 _1588_ (.B(_0806_),
    .C(_0793_),
    .A(_0787_),
    .Y(_0815_),
    .D(_0808_));
 sg13g2_a21oi_1 _1589_ (.A1(_0814_),
    .A2(_0815_),
    .Y(_0816_),
    .B1(net17));
 sg13g2_xor2_1 _1590_ (.B(_0816_),
    .A(\top_inst.sprite_movement_inst.sprite_y[6] ),
    .X(_0155_));
 sg13g2_nor4_1 _1591_ (.A(_0806_),
    .B(\top_inst.sprite_movement_inst.sprite_y[6] ),
    .C(_0793_),
    .D(_0810_),
    .Y(_0817_));
 sg13g2_and4_1 _1592_ (.A(_0806_),
    .B(\top_inst.sprite_movement_inst.sprite_y[6] ),
    .C(_0793_),
    .D(_0810_),
    .X(_0818_));
 sg13g2_nor2_1 _1593_ (.A(_0817_),
    .B(_0818_),
    .Y(_0819_));
 sg13g2_nor2_1 _1594_ (.A(_0743_),
    .B(_0819_),
    .Y(_0820_));
 sg13g2_xor2_1 _1595_ (.B(_0820_),
    .A(\top_inst.sprite_movement_inst.sprite_y[7] ),
    .X(_0156_));
 sg13g2_or2_1 _1596_ (.X(_0821_),
    .B(\top_inst.sprite_movement_inst.sprite_y[6] ),
    .A(\top_inst.sprite_movement_inst.sprite_y[7] ));
 sg13g2_nand2_1 _1597_ (.Y(_0822_),
    .A(_0786_),
    .B(_0813_));
 sg13g2_nor3_1 _1598_ (.A(net16),
    .B(_0821_),
    .C(_0822_),
    .Y(_0823_));
 sg13g2_nand4_1 _1599_ (.B(_0791_),
    .C(_0802_),
    .A(_0798_),
    .Y(_0824_),
    .D(_0806_));
 sg13g2_nor4_1 _1600_ (.A(_0786_),
    .B(_0743_),
    .C(_0821_),
    .D(_0824_),
    .Y(_0825_));
 sg13g2_o21ai_1 _1601_ (.B1(_0787_),
    .Y(_0826_),
    .A1(_0788_),
    .A2(_0825_));
 sg13g2_o21ai_1 _1602_ (.B1(_0826_),
    .Y(_0157_),
    .A1(_0793_),
    .A2(_0823_));
 sg13g2_nand3_1 _1603_ (.B(_0559_),
    .C(_0586_),
    .A(_0565_),
    .Y(_0827_));
 sg13g2_nand4_1 _1604_ (.B(net43),
    .C(_0553_),
    .A(_0583_),
    .Y(_0828_),
    .D(\top_inst.background_inst.cur_time[7] ));
 sg13g2_nor2_1 _1605_ (.A(_0827_),
    .B(_0828_),
    .Y(_0829_));
 sg13g2_nand2_1 _1606_ (.Y(_0830_),
    .A(next_frame),
    .B(_0829_));
 sg13g2_or2_1 _1607_ (.X(_0831_),
    .B(_0571_),
    .A(net40));
 sg13g2_or4_1 _1608_ (.A(_0565_),
    .B(net43),
    .C(_0553_),
    .D(\top_inst.background_inst.cur_time[7] ),
    .X(_0832_));
 sg13g2_nor4_1 _1609_ (.A(_0583_),
    .B(_0567_),
    .C(_0831_),
    .D(_0832_),
    .Y(_0833_));
 sg13g2_a22oi_1 _1610_ (.Y(_0174_),
    .B1(_0833_),
    .B2(next_frame),
    .A2(_0830_),
    .A1(_0560_));
 sg13g2_buf_1 _1611_ (.A(_0491_),
    .X(_0834_));
 sg13g2_or3_1 _1612_ (.A(\top_inst.spi_receiver_inst.registers[4][0] ),
    .B(\top_inst.spi_receiver_inst.registers[4][2] ),
    .C(\top_inst.spi_receiver_inst.registers[4][1] ),
    .X(_0835_));
 sg13g2_nand3_1 _1613_ (.B(\top_inst.spi_receiver_inst.registers[4][3] ),
    .C(_0835_),
    .A(\top_inst.spi_receiver_inst.registers[4][4] ),
    .Y(_0836_));
 sg13g2_buf_1 _1614_ (.A(\top_inst.misc[2] ),
    .X(_0837_));
 sg13g2_nor3_1 _1615_ (.A(net28),
    .B(\top_inst.spi_receiver_inst.registers[4][7] ),
    .C(\top_inst.spi_receiver_inst.registers[4][5] ),
    .Y(_0838_));
 sg13g2_nand3b_1 _1616_ (.B(net37),
    .C(_0756_),
    .Y(_0839_),
    .A_N(_0758_));
 sg13g2_nand2b_1 _1617_ (.Y(_0840_),
    .B(\top_inst.misc[2] ),
    .A_N(\top_inst.sprite_movement_inst.sprite_x[7] ));
 sg13g2_nor2_1 _1618_ (.A(_0766_),
    .B(_0840_),
    .Y(_0841_));
 sg13g2_or3_1 _1619_ (.A(\top_inst.misc[2] ),
    .B(\top_inst.spi_receiver_inst.registers[4][7] ),
    .C(\top_inst.spi_receiver_inst.registers[4][6] ),
    .X(_0842_));
 sg13g2_o21ai_1 _1620_ (.B1(_0842_),
    .Y(_0843_),
    .A1(_0773_),
    .A2(_0840_));
 sg13g2_a221oi_1 _1621_ (.B2(_0841_),
    .C1(_0843_),
    .B1(_0839_),
    .A1(_0836_),
    .Y(_0844_),
    .A2(_0838_));
 sg13g2_buf_1 _1622_ (.A(_0844_),
    .X(_0845_));
 sg13g2_buf_1 _1623_ (.A(net28),
    .X(_0846_));
 sg13g2_nor2b_1 _1624_ (.A(net28),
    .B_N(\top_inst.spi_receiver_inst.registers[4][0] ),
    .Y(_0847_));
 sg13g2_a21oi_1 _1625_ (.A1(net27),
    .A2(_0741_),
    .Y(_0848_),
    .B1(_0847_));
 sg13g2_nor3_1 _1626_ (.A(_0491_),
    .B(_0845_),
    .C(_0848_),
    .Y(_0849_));
 sg13g2_a21o_1 _1627_ (.A2(net25),
    .A1(\top_inst.sprite_x[0] ),
    .B1(_0849_),
    .X(_0158_));
 sg13g2_nor2b_1 _1628_ (.A(net28),
    .B_N(\top_inst.spi_receiver_inst.registers[4][1] ),
    .Y(_0850_));
 sg13g2_a21oi_1 _1629_ (.A1(net27),
    .A2(_0745_),
    .Y(_0851_),
    .B1(_0850_));
 sg13g2_nor3_1 _1630_ (.A(_0491_),
    .B(_0845_),
    .C(_0851_),
    .Y(_0852_));
 sg13g2_a21o_1 _1631_ (.A2(net25),
    .A1(\top_inst.sprite_x[1] ),
    .B1(_0852_),
    .X(_0159_));
 sg13g2_nor2b_1 _1632_ (.A(net28),
    .B_N(\top_inst.spi_receiver_inst.registers[4][2] ),
    .Y(_0853_));
 sg13g2_a21oi_1 _1633_ (.A1(net27),
    .A2(_0750_),
    .Y(_0854_),
    .B1(_0853_));
 sg13g2_nor3_1 _1634_ (.A(_0491_),
    .B(_0845_),
    .C(_0854_),
    .Y(_0855_));
 sg13g2_a21o_1 _1635_ (.A2(net25),
    .A1(_0600_),
    .B1(_0855_),
    .X(_0160_));
 sg13g2_inv_1 _1636_ (.Y(_0856_),
    .A(_0599_));
 sg13g2_mux2_1 _1637_ (.A0(\top_inst.spi_receiver_inst.registers[4][3] ),
    .A1(_0756_),
    .S(net27),
    .X(_0857_));
 sg13g2_buf_1 _1638_ (.A(net24),
    .X(_0858_));
 sg13g2_o21ai_1 _1639_ (.B1(net21),
    .Y(_0859_),
    .A1(_0845_),
    .A2(_0857_));
 sg13g2_o21ai_1 _1640_ (.B1(_0859_),
    .Y(_0161_),
    .A1(_0856_),
    .A2(net22));
 sg13g2_inv_1 _1641_ (.Y(_0860_),
    .A(\top_inst.sprite_x[4] ));
 sg13g2_mux2_1 _1642_ (.A0(\top_inst.spi_receiver_inst.registers[4][4] ),
    .A1(_0762_),
    .S(net27),
    .X(_0861_));
 sg13g2_o21ai_1 _1643_ (.B1(net21),
    .Y(_0862_),
    .A1(_0845_),
    .A2(_0861_));
 sg13g2_o21ai_1 _1644_ (.B1(_0862_),
    .Y(_0162_),
    .A1(_0860_),
    .A2(net22));
 sg13g2_mux2_1 _1645_ (.A0(\top_inst.spi_receiver_inst.registers[4][5] ),
    .A1(_0766_),
    .S(net27),
    .X(_0863_));
 sg13g2_nand3_1 _1646_ (.B(_0843_),
    .C(_0863_),
    .A(net24),
    .Y(_0864_));
 sg13g2_o21ai_1 _1647_ (.B1(_0864_),
    .Y(_0163_),
    .A1(_0607_),
    .A2(net22));
 sg13g2_nand2_1 _1648_ (.Y(_0865_),
    .A(\top_inst.sprite_x[6] ),
    .B(net25));
 sg13g2_o21ai_1 _1649_ (.B1(_0865_),
    .Y(_0164_),
    .A1(net25),
    .A2(_0843_));
 sg13g2_nor2_1 _1650_ (.A(_0635_),
    .B(net23),
    .Y(_0165_));
 sg13g2_inv_1 _1651_ (.Y(_0866_),
    .A(\top_inst.sprite_y[0] ));
 sg13g2_nor2_1 _1652_ (.A(\top_inst.sprite_movement_inst.sprite_y[7] ),
    .B(\top_inst.sprite_movement_inst.sprite_y[6] ),
    .Y(_0867_));
 sg13g2_nor3_1 _1653_ (.A(_0837_),
    .B(\top_inst.spi_receiver_inst.registers[5][7] ),
    .C(\top_inst.spi_receiver_inst.registers[5][6] ),
    .Y(_0868_));
 sg13g2_a21oi_2 _1654_ (.B1(_0868_),
    .Y(_0869_),
    .A2(_0867_),
    .A1(net28));
 sg13g2_mux2_1 _1655_ (.A0(\top_inst.spi_receiver_inst.registers[5][0] ),
    .A1(_0786_),
    .S(net27),
    .X(_0870_));
 sg13g2_o21ai_1 _1656_ (.B1(net21),
    .Y(_0871_),
    .A1(_0869_),
    .A2(_0870_));
 sg13g2_o21ai_1 _1657_ (.B1(_0871_),
    .Y(_0166_),
    .A1(_0866_),
    .A2(net22));
 sg13g2_inv_1 _1658_ (.Y(_0872_),
    .A(\top_inst.sprite_y[1] ));
 sg13g2_mux2_1 _1659_ (.A0(\top_inst.spi_receiver_inst.registers[5][1] ),
    .A1(_0787_),
    .S(_0846_),
    .X(_0873_));
 sg13g2_o21ai_1 _1660_ (.B1(net21),
    .Y(_0874_),
    .A1(_0869_),
    .A2(_0873_));
 sg13g2_o21ai_1 _1661_ (.B1(_0874_),
    .Y(_0167_),
    .A1(_0872_),
    .A2(net22));
 sg13g2_nor2_1 _1662_ (.A(_0846_),
    .B(\top_inst.spi_receiver_inst.registers[5][2] ),
    .Y(_0875_));
 sg13g2_a21oi_1 _1663_ (.A1(net27),
    .A2(_0792_),
    .Y(_0876_),
    .B1(_0875_));
 sg13g2_o21ai_1 _1664_ (.B1(net21),
    .Y(_0877_),
    .A1(_0869_),
    .A2(_0876_));
 sg13g2_o21ai_1 _1665_ (.B1(_0877_),
    .Y(_0168_),
    .A1(_0723_),
    .A2(net21));
 sg13g2_mux2_1 _1666_ (.A0(\top_inst.spi_receiver_inst.registers[5][3] ),
    .A1(_0798_),
    .S(_0837_),
    .X(_0878_));
 sg13g2_o21ai_1 _1667_ (.B1(net24),
    .Y(_0879_),
    .A1(_0869_),
    .A2(_0878_));
 sg13g2_o21ai_1 _1668_ (.B1(_0879_),
    .Y(_0169_),
    .A1(_0717_),
    .A2(_0858_));
 sg13g2_inv_1 _1669_ (.Y(_0880_),
    .A(_0646_));
 sg13g2_mux2_1 _1670_ (.A0(\top_inst.spi_receiver_inst.registers[5][4] ),
    .A1(_0802_),
    .S(net28),
    .X(_0881_));
 sg13g2_o21ai_1 _1671_ (.B1(net24),
    .Y(_0882_),
    .A1(_0869_),
    .A2(_0881_));
 sg13g2_o21ai_1 _1672_ (.B1(_0882_),
    .Y(_0170_),
    .A1(_0880_),
    .A2(net21));
 sg13g2_mux2_1 _1673_ (.A0(\top_inst.spi_receiver_inst.registers[5][5] ),
    .A1(_0806_),
    .S(net28),
    .X(_0883_));
 sg13g2_o21ai_1 _1674_ (.B1(net24),
    .Y(_0884_),
    .A1(_0869_),
    .A2(_0883_));
 sg13g2_o21ai_1 _1675_ (.B1(_0884_),
    .Y(_0171_),
    .A1(_0643_),
    .A2(net21));
 sg13g2_nor2_1 _1676_ (.A(_0641_),
    .B(net23),
    .Y(_0172_));
 sg13g2_nor2_1 _1677_ (.A(_0672_),
    .B(net23),
    .Y(_0173_));
 sg13g2_nand2b_1 _1678_ (.Y(_0885_),
    .B(_0492_),
    .A_N(_0513_));
 sg13g2_buf_1 _1679_ (.A(_0885_),
    .X(_0886_));
 sg13g2_inv_1 _1680_ (.Y(_0887_),
    .A(net20));
 sg13g2_a22oi_1 _1681_ (.Y(_0888_),
    .B1(_0887_),
    .B2(_0042_),
    .A2(_0491_),
    .A1(net32));
 sg13g2_inv_1 _1682_ (.Y(_0175_),
    .A(_0888_));
 sg13g2_buf_1 _1683_ (.A(_0502_),
    .X(_0889_));
 sg13g2_and2_1 _1684_ (.A(net35),
    .B(_0501_),
    .X(_0890_));
 sg13g2_buf_1 _1685_ (.A(_0890_),
    .X(_0891_));
 sg13g2_nand3_1 _1686_ (.B(net30),
    .C(_0891_),
    .A(net36),
    .Y(_0892_));
 sg13g2_or2_1 _1687_ (.X(_0893_),
    .B(_0892_),
    .A(_0722_));
 sg13g2_nor2_1 _1688_ (.A(_0662_),
    .B(_0893_),
    .Y(_0894_));
 sg13g2_nand3_1 _1689_ (.B(_0509_),
    .C(_0894_),
    .A(_0660_),
    .Y(_0895_));
 sg13g2_a21oi_1 _1690_ (.A1(_0510_),
    .A2(_0895_),
    .Y(_0896_),
    .B1(net20));
 sg13g2_a21o_1 _1691_ (.A2(net25),
    .A1(_0048_),
    .B1(_0896_),
    .X(_0176_));
 sg13g2_inv_1 _1692_ (.Y(_0897_),
    .A(net47));
 sg13g2_nand2_1 _1693_ (.Y(_0898_),
    .A(_0897_),
    .B(net32));
 sg13g2_o21ai_1 _1694_ (.B1(net24),
    .Y(_0899_),
    .A1(net32),
    .A2(_0513_));
 sg13g2_nand2_1 _1695_ (.Y(_0900_),
    .A(net47),
    .B(_0899_));
 sg13g2_o21ai_1 _1696_ (.B1(_0900_),
    .Y(_0177_),
    .A1(net20),
    .A2(_0898_));
 sg13g2_inv_1 _1697_ (.Y(_0901_),
    .A(_0049_));
 sg13g2_a21oi_1 _1698_ (.A1(net47),
    .A2(net32),
    .Y(_0902_),
    .B1(net31));
 sg13g2_o21ai_1 _1699_ (.B1(_0887_),
    .Y(_0903_),
    .A1(_0501_),
    .A2(_0902_));
 sg13g2_o21ai_1 _1700_ (.B1(_0903_),
    .Y(_0178_),
    .A1(_0901_),
    .A2(_0858_));
 sg13g2_xor2_1 _1701_ (.B(_0501_),
    .A(_0039_),
    .X(_0904_));
 sg13g2_nand2_1 _1702_ (.Y(_0905_),
    .A(net35),
    .B(_0834_));
 sg13g2_o21ai_1 _1703_ (.B1(_0905_),
    .Y(_0179_),
    .A1(net20),
    .A2(_0904_));
 sg13g2_nand2_1 _1704_ (.Y(_0906_),
    .A(_0887_),
    .B(_0891_));
 sg13g2_o21ai_1 _1705_ (.B1(_0523_),
    .Y(_0907_),
    .A1(_0513_),
    .A2(_0891_));
 sg13g2_nand2_1 _1706_ (.Y(_0908_),
    .A(net30),
    .B(_0907_));
 sg13g2_o21ai_1 _1707_ (.B1(_0908_),
    .Y(_0180_),
    .A1(net30),
    .A2(_0906_));
 sg13g2_a21o_1 _1708_ (.A2(_0891_),
    .A1(net30),
    .B1(net36),
    .X(_0909_));
 sg13g2_and2_1 _1709_ (.A(_0892_),
    .B(_0909_),
    .X(_0910_));
 sg13g2_nand2_1 _1710_ (.Y(_0911_),
    .A(_0050_),
    .B(_0834_));
 sg13g2_o21ai_1 _1711_ (.B1(_0911_),
    .Y(_0181_),
    .A1(_0886_),
    .A2(_0910_));
 sg13g2_xnor2_1 _1712_ (.Y(_0912_),
    .A(net46),
    .B(_0892_));
 sg13g2_nand2_1 _1713_ (.Y(_0913_),
    .A(_0051_),
    .B(net25));
 sg13g2_o21ai_1 _1714_ (.B1(_0913_),
    .Y(_0182_),
    .A1(net20),
    .A2(_0912_));
 sg13g2_xnor2_1 _1715_ (.Y(_0914_),
    .A(_0507_),
    .B(_0893_));
 sg13g2_nand2_1 _1716_ (.Y(_0915_),
    .A(_0052_),
    .B(net25));
 sg13g2_o21ai_1 _1717_ (.B1(_0915_),
    .Y(_0183_),
    .A1(net20),
    .A2(_0914_));
 sg13g2_xor2_1 _1718_ (.B(_0894_),
    .A(_0660_),
    .X(_0916_));
 sg13g2_nand2_1 _1719_ (.Y(_0917_),
    .A(_0053_),
    .B(_0491_));
 sg13g2_o21ai_1 _1720_ (.B1(_0917_),
    .Y(_0184_),
    .A1(net20),
    .A2(_0916_));
 sg13g2_nand2_1 _1721_ (.Y(_0918_),
    .A(net39),
    .B(_0894_));
 sg13g2_xnor2_1 _1722_ (.Y(_0919_),
    .A(_0509_),
    .B(_0918_));
 sg13g2_nand2_1 _1723_ (.Y(_0920_),
    .A(_0054_),
    .B(_0491_));
 sg13g2_o21ai_1 _1724_ (.B1(_0920_),
    .Y(_0185_),
    .A1(net20),
    .A2(_0919_));
 sg13g2_inv_1 _1725_ (.Y(_0055_),
    .A(\top_inst.sprite_data_inst.sprite_data[103] ));
 sg13g2_inv_1 _1726_ (.Y(_0056_),
    .A(\top_inst.sprite_data_inst.sprite_data[115] ));
 sg13g2_inv_1 _1727_ (.Y(_0057_),
    .A(\top_inst.sprite_data_inst.sprite_data[127] ));
 sg13g2_inv_1 _1728_ (.Y(_0058_),
    .A(\top_inst.sprite_data_inst.sprite_data[136] ));
 sg13g2_inv_1 _1729_ (.Y(_0059_),
    .A(\top_inst.sprite_data_inst.sprite_data[137] ));
 sg13g2_inv_1 _1730_ (.Y(_0060_),
    .A(\top_inst.sprite_data_inst.sprite_data[138] ));
 sg13g2_inv_1 _1731_ (.Y(_0061_),
    .A(\top_inst.sprite_data_inst.sprite_data[139] ));
 sg13g2_inv_1 _1732_ (.Y(_0062_),
    .A(\top_inst.sprite_data_inst.sprite_data[26] ));
 sg13g2_inv_1 _1733_ (.Y(_0063_),
    .A(\top_inst.sprite_data_inst.sprite_data[27] ));
 sg13g2_inv_1 _1734_ (.Y(_0064_),
    .A(\top_inst.sprite_data_inst.sprite_data[28] ));
 sg13g2_inv_1 _1735_ (.Y(_0065_),
    .A(\top_inst.sprite_data_inst.sprite_data[29] ));
 sg13g2_inv_1 _1736_ (.Y(_0066_),
    .A(\top_inst.sprite_data_inst.sprite_data[30] ));
 sg13g2_inv_1 _1737_ (.Y(_0067_),
    .A(\top_inst.sprite_data_inst.sprite_data[37] ));
 sg13g2_inv_1 _1738_ (.Y(_0068_),
    .A(\top_inst.sprite_data_inst.sprite_data[38] ));
 sg13g2_inv_1 _1739_ (.Y(_0069_),
    .A(\top_inst.sprite_data_inst.sprite_data[39] ));
 sg13g2_inv_1 _1740_ (.Y(_0070_),
    .A(\top_inst.sprite_data_inst.sprite_data[40] ));
 sg13g2_inv_1 _1741_ (.Y(_0071_),
    .A(\top_inst.sprite_data_inst.sprite_data[4] ));
 sg13g2_inv_1 _1742_ (.Y(_0072_),
    .A(\top_inst.sprite_data_inst.sprite_data[41] ));
 sg13g2_inv_1 _1743_ (.Y(_0073_),
    .A(\top_inst.sprite_data_inst.sprite_data[42] ));
 sg13g2_inv_1 _1744_ (.Y(_0074_),
    .A(\top_inst.sprite_data_inst.sprite_data[5] ));
 sg13g2_inv_1 _1745_ (.Y(_0075_),
    .A(\top_inst.sprite_data_inst.sprite_data[52] ));
 sg13g2_inv_1 _1746_ (.Y(_0076_),
    .A(\top_inst.sprite_data_inst.sprite_data[60] ));
 sg13g2_inv_1 _1747_ (.Y(_0077_),
    .A(\top_inst.sprite_data_inst.sprite_data[6] ));
 sg13g2_inv_1 _1748_ (.Y(_0078_),
    .A(\top_inst.sprite_data_inst.sprite_data[64] ));
 sg13g2_inv_1 _1749_ (.Y(_0079_),
    .A(\top_inst.sprite_data_inst.sprite_data[65] ));
 sg13g2_inv_1 _1750_ (.Y(_0080_),
    .A(\top_inst.sprite_data_inst.sprite_data[66] ));
 sg13g2_inv_1 _1751_ (.Y(_0081_),
    .A(\top_inst.sprite_data_inst.sprite_data[67] ));
 sg13g2_inv_1 _1752_ (.Y(_0082_),
    .A(\top_inst.sprite_data_inst.sprite_data[68] ));
 sg13g2_inv_1 _1753_ (.Y(_0083_),
    .A(\top_inst.sprite_data_inst.sprite_data[69] ));
 sg13g2_inv_1 _1754_ (.Y(_0084_),
    .A(\top_inst.sprite_data_inst.sprite_data[7] ));
 sg13g2_inv_1 _1755_ (.Y(_0085_),
    .A(\top_inst.sprite_data_inst.sprite_data[72] ));
 sg13g2_inv_1 _1756_ (.Y(_0086_),
    .A(\top_inst.sprite_data_inst.sprite_data[76] ));
 sg13g2_inv_1 _1757_ (.Y(_0087_),
    .A(\top_inst.sprite_data_inst.sprite_data[77] ));
 sg13g2_inv_1 _1758_ (.Y(_0088_),
    .A(\top_inst.sprite_data_inst.sprite_data[78] ));
 sg13g2_inv_1 _1759_ (.Y(_0089_),
    .A(\top_inst.sprite_data_inst.sprite_data[79] ));
 sg13g2_inv_1 _1760_ (.Y(_0090_),
    .A(\top_inst.sprite_data_inst.sprite_data[80] ));
 sg13g2_inv_1 _1761_ (.Y(_0091_),
    .A(\top_inst.sprite_data_inst.sprite_data[8] ));
 sg13g2_inv_1 _1762_ (.Y(_0092_),
    .A(\top_inst.sprite_data_inst.sprite_data[81] ));
 sg13g2_inv_1 _1763_ (.Y(_0093_),
    .A(\top_inst.sprite_data_inst.sprite_data[84] ));
 sg13g2_inv_1 _1764_ (.Y(_0094_),
    .A(\top_inst.sprite_data_inst.sprite_data[88] ));
 sg13g2_inv_1 _1765_ (.Y(_0095_),
    .A(\top_inst.sprite_data_inst.sprite_data[91] ));
 sg13g2_inv_1 _1766_ (.Y(_0096_),
    .A(\top_inst.sprite_data_inst.sprite_data[96] ));
 sg13g2_inv_1 _1767_ (.Y(_0097_),
    .A(\top_inst.sprite_data_inst.sprite_data[100] ));
 sg13g2_nor2_1 _1768_ (.A(_0537_),
    .B(_0538_),
    .Y(_0186_));
 sg13g2_nand2_1 _1769_ (.Y(_0187_),
    .A(_0474_),
    .B(_0186_));
 sg13g2_xnor2_1 _1770_ (.Y(_0188_),
    .A(net48),
    .B(_0187_));
 sg13g2_nor2_1 _1771_ (.A(net22),
    .B(_0188_),
    .Y(_0098_));
 sg13g2_nand2_1 _1772_ (.Y(_0189_),
    .A(\top_inst.background_inst.counter_h[8] ),
    .B(_0186_));
 sg13g2_nand3_1 _1773_ (.B(_0472_),
    .C(net51),
    .A(net48),
    .Y(_0190_));
 sg13g2_nand2b_1 _1774_ (.Y(_0191_),
    .B(_0489_),
    .A_N(_0472_));
 sg13g2_o21ai_1 _1775_ (.B1(_0191_),
    .Y(_0099_),
    .A1(_0189_),
    .A2(_0190_));
 sg13g2_o21ai_1 _1776_ (.B1(_0606_),
    .Y(_0192_),
    .A1(_0537_),
    .A2(_0538_));
 sg13g2_a21oi_1 _1777_ (.A1(_0189_),
    .A2(_0192_),
    .Y(_0100_),
    .B1(_0534_));
 sg13g2_nand2b_1 _1778_ (.Y(_0193_),
    .B(_0189_),
    .A_N(net51));
 sg13g2_a21oi_1 _1779_ (.A1(_0187_),
    .A2(_0193_),
    .Y(_0101_),
    .B1(_0534_));
 sg13g2_nand3_1 _1780_ (.B(_0472_),
    .C(_0474_),
    .A(_0488_),
    .Y(_0194_));
 sg13g2_nor3_1 _1781_ (.A(_0478_),
    .B(_0479_),
    .C(_0480_),
    .Y(_0195_));
 sg13g2_nand3_1 _1782_ (.B(_0477_),
    .C(_0195_),
    .A(_0475_),
    .Y(_0196_));
 sg13g2_inv_1 _1783_ (.Y(_0197_),
    .A(\top_inst.background_inst.counter_h[5] ));
 sg13g2_nor3_1 _1784_ (.A(net45),
    .B(_0197_),
    .C(_0476_),
    .Y(_0198_));
 sg13g2_a21oi_1 _1785_ (.A1(_0038_),
    .A2(_0196_),
    .Y(_0199_),
    .B1(_0198_));
 sg13g2_nor2_1 _1786_ (.A(_0484_),
    .B(_0199_),
    .Y(_0200_));
 sg13g2_xnor2_1 _1787_ (.Y(_0201_),
    .A(_0537_),
    .B(_0200_));
 sg13g2_nor2_1 _1788_ (.A(_0194_),
    .B(_0201_),
    .Y(hsync));
 sg13g2_mux2_1 _1789_ (.A0(\top_inst.sprite_access_inst.sprite_data ),
    .A1(net167),
    .S(net2),
    .X(\top_inst.sprite_data_inst.new_sprite_data ));
 sg13g2_a22oi_1 _1790_ (.Y(_0202_),
    .B1(net18),
    .B2(_0736_),
    .A2(_0544_),
    .A1(net2));
 sg13g2_inv_1 _1791_ (.Y(\top_inst.sprite_data_inst.shiftf ),
    .A(_0202_));
 sg13g2_and3_1 _1792_ (.X(_0203_),
    .A(net46),
    .B(_0507_),
    .C(net36));
 sg13g2_nand4_1 _1793_ (.B(_0509_),
    .C(_0510_),
    .A(net39),
    .Y(_0204_),
    .D(_0203_));
 sg13g2_nor3_1 _1794_ (.A(net47),
    .B(net32),
    .C(net35),
    .Y(_0205_));
 sg13g2_inv_1 _1795_ (.Y(_0206_),
    .A(_0495_));
 sg13g2_nor2b_1 _1796_ (.A(net30),
    .B_N(net32),
    .Y(_0207_));
 sg13g2_o21ai_1 _1797_ (.B1(_0203_),
    .Y(_0208_),
    .A1(net31),
    .A2(_0207_));
 sg13g2_nor2_1 _1798_ (.A(net47),
    .B(_0206_),
    .Y(_0209_));
 sg13g2_a22oi_1 _1799_ (.Y(_0210_),
    .B1(_0208_),
    .B2(_0209_),
    .A2(_0206_),
    .A1(net31));
 sg13g2_nor4_1 _1800_ (.A(net30),
    .B(_0204_),
    .C(_0205_),
    .D(_0210_),
    .Y(\top_inst.timing_ver.sync ));
 sg13g2_inv_1 _1801_ (.Y(_0211_),
    .A(\top_inst.background_inst.bg_select[1] ));
 sg13g2_buf_2 _1802_ (.A(\top_inst.misc[3] ),
    .X(_0212_));
 sg13g2_nor2_1 _1803_ (.A(_0212_),
    .B(_0737_),
    .Y(_0213_));
 sg13g2_nand3_1 _1804_ (.B(net32),
    .C(_0042_),
    .A(_0897_),
    .Y(_0214_));
 sg13g2_or2_1 _1805_ (.X(_0215_),
    .B(_0889_),
    .A(net35));
 sg13g2_a21oi_1 _1806_ (.A1(net31),
    .A2(_0214_),
    .Y(_0216_),
    .B1(_0215_));
 sg13g2_or2_1 _1807_ (.X(_0217_),
    .B(_0216_),
    .A(_0204_));
 sg13g2_and2_1 _1808_ (.A(_0194_),
    .B(_0217_),
    .X(_0218_));
 sg13g2_o21ai_1 _1809_ (.B1(_0218_),
    .Y(_0219_),
    .A1(_0731_),
    .A2(_0213_));
 sg13g2_or2_1 _1810_ (.X(_0220_),
    .B(_0219_),
    .A(_0211_));
 sg13g2_inv_1 _1811_ (.Y(_0221_),
    .A(\top_inst.background_inst.color1[5] ));
 sg13g2_inv_1 _1812_ (.Y(_0222_),
    .A(\top_inst.background_inst.color3[5] ));
 sg13g2_inv_1 _1813_ (.Y(_0223_),
    .A(\top_inst.background_inst.color2[5] ));
 sg13g2_inv_1 _1814_ (.Y(_0224_),
    .A(\top_inst.background_inst.color4[5] ));
 sg13g2_xnor2_1 _1815_ (.Y(_0225_),
    .A(_0505_),
    .B(_0583_));
 sg13g2_nor2b_1 _1816_ (.A(_0225_),
    .B_N(\top_inst.background_inst.bg_select[0] ),
    .Y(_0226_));
 sg13g2_and2_1 _1817_ (.A(\top_inst.background_inst.bg_select[0] ),
    .B(_0225_),
    .X(_0227_));
 sg13g2_nor2_2 _1818_ (.A(\top_inst.background_inst.counter_v[1] ),
    .B(_0555_),
    .Y(_0228_));
 sg13g2_nor2_1 _1819_ (.A(_0499_),
    .B(net43),
    .Y(_0229_));
 sg13g2_nand2_1 _1820_ (.Y(_0230_),
    .A(_0498_),
    .B(_0552_));
 sg13g2_a221oi_1 _1821_ (.B2(_0498_),
    .C1(net42),
    .B1(_0552_),
    .A1(_0497_),
    .Y(_0231_),
    .A2(net43));
 sg13g2_a221oi_1 _1822_ (.B2(_0230_),
    .C1(_0231_),
    .B1(_0229_),
    .A1(_0566_),
    .Y(_0232_),
    .A2(_0228_));
 sg13g2_inv_1 _1823_ (.Y(_0233_),
    .A(_0499_));
 sg13g2_nor2_1 _1824_ (.A(net47),
    .B(net31),
    .Y(_0234_));
 sg13g2_nor2_1 _1825_ (.A(_0499_),
    .B(\top_inst.background_inst.cur_time[2] ),
    .Y(_0235_));
 sg13g2_a221oi_1 _1826_ (.B2(_0230_),
    .C1(_0235_),
    .B1(_0234_),
    .A1(_0233_),
    .Y(_0236_),
    .A2(_0228_));
 sg13g2_inv_1 _1827_ (.Y(_0237_),
    .A(\top_inst.background_inst.cur_time[3] ));
 sg13g2_nor2_1 _1828_ (.A(_0206_),
    .B(_0237_),
    .Y(_0238_));
 sg13g2_a21o_1 _1829_ (.A2(_0236_),
    .A1(_0232_),
    .B1(_0238_),
    .X(_0239_));
 sg13g2_buf_1 _1830_ (.A(_0237_),
    .X(_0240_));
 sg13g2_nand2_1 _1831_ (.Y(_0241_),
    .A(_0206_),
    .B(net29));
 sg13g2_and2_1 _1832_ (.A(_0493_),
    .B(net40),
    .X(_0242_));
 sg13g2_a221oi_1 _1833_ (.B2(_0241_),
    .C1(_0242_),
    .B1(_0239_),
    .A1(net30),
    .Y(_0243_),
    .A2(_0571_));
 sg13g2_nor2_1 _1834_ (.A(net30),
    .B(_0571_),
    .Y(_0244_));
 sg13g2_nand2_1 _1835_ (.Y(_0245_),
    .A(_0493_),
    .B(net40));
 sg13g2_nor2_1 _1836_ (.A(_0493_),
    .B(net40),
    .Y(_0246_));
 sg13g2_a21oi_1 _1837_ (.A1(_0244_),
    .A2(_0245_),
    .Y(_0247_),
    .B1(_0246_));
 sg13g2_nand2b_1 _1838_ (.Y(_0248_),
    .B(_0247_),
    .A_N(_0243_));
 sg13g2_mux2_1 _1839_ (.A0(_0226_),
    .A1(_0227_),
    .S(_0248_),
    .X(_0249_));
 sg13g2_buf_1 _1840_ (.A(_0249_),
    .X(_0250_));
 sg13g2_a21oi_1 _1841_ (.A1(_0499_),
    .A2(\top_inst.background_inst.cur_time[2] ),
    .Y(_0251_),
    .B1(_0478_));
 sg13g2_nor2_1 _1842_ (.A(_0235_),
    .B(_0251_),
    .Y(_0252_));
 sg13g2_xnor2_1 _1843_ (.Y(_0253_),
    .A(\top_inst.background_inst.cur_time[3] ),
    .B(_0252_));
 sg13g2_nand2_1 _1844_ (.Y(_0254_),
    .A(net45),
    .B(net35));
 sg13g2_or2_1 _1845_ (.X(_0255_),
    .B(net35),
    .A(net45));
 sg13g2_xnor2_1 _1846_ (.Y(_0256_),
    .A(_0476_),
    .B(_0502_));
 sg13g2_xnor2_1 _1847_ (.Y(_0257_),
    .A(_0571_),
    .B(_0256_));
 sg13g2_mux2_1 _1848_ (.A0(_0254_),
    .A1(_0255_),
    .S(_0257_),
    .X(_0258_));
 sg13g2_xor2_1 _1849_ (.B(_0495_),
    .A(net45),
    .X(_0259_));
 sg13g2_nand2_1 _1850_ (.Y(_0260_),
    .A(net31),
    .B(net42));
 sg13g2_o21ai_1 _1851_ (.B1(_0478_),
    .Y(_0261_),
    .A1(_0499_),
    .A2(net42));
 sg13g2_nand4_1 _1852_ (.B(_0259_),
    .C(_0260_),
    .A(net29),
    .Y(_0262_),
    .D(_0261_));
 sg13g2_xnor2_1 _1853_ (.Y(_0263_),
    .A(net45),
    .B(_0495_));
 sg13g2_or4_1 _1854_ (.A(_0237_),
    .B(_0263_),
    .C(_0235_),
    .D(_0251_),
    .X(_0264_));
 sg13g2_xor2_1 _1855_ (.B(_0256_),
    .A(_0571_),
    .X(_0265_));
 sg13g2_mux2_1 _1856_ (.A0(_0262_),
    .A1(_0264_),
    .S(_0265_),
    .X(_0266_));
 sg13g2_o21ai_1 _1857_ (.B1(_0266_),
    .Y(_0267_),
    .A1(_0253_),
    .A2(_0258_));
 sg13g2_xnor2_1 _1858_ (.Y(_0268_),
    .A(net49),
    .B(_0225_));
 sg13g2_a21oi_1 _1859_ (.A1(_0197_),
    .A2(_0245_),
    .Y(_0269_),
    .B1(_0246_));
 sg13g2_xnor2_1 _1860_ (.Y(_0270_),
    .A(_0268_),
    .B(_0269_));
 sg13g2_nand2_2 _1861_ (.Y(_0271_),
    .A(_0502_),
    .B(_0571_));
 sg13g2_o21ai_1 _1862_ (.B1(_0476_),
    .Y(_0272_),
    .A1(_0502_),
    .A2(_0571_));
 sg13g2_nand2_1 _1863_ (.Y(_0273_),
    .A(_0271_),
    .B(_0272_));
 sg13g2_xnor2_1 _1864_ (.Y(_0274_),
    .A(_0493_),
    .B(net40));
 sg13g2_xnor2_1 _1865_ (.Y(_0275_),
    .A(net50),
    .B(_0274_));
 sg13g2_xnor2_1 _1866_ (.Y(_0276_),
    .A(_0273_),
    .B(_0275_));
 sg13g2_nor2_1 _1867_ (.A(_0270_),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_o21ai_1 _1868_ (.B1(_0498_),
    .Y(_0278_),
    .A1(_0480_),
    .A2(_0552_));
 sg13g2_nand2_1 _1869_ (.Y(_0279_),
    .A(_0480_),
    .B(_0552_));
 sg13g2_xor2_1 _1870_ (.B(\top_inst.background_inst.cur_time[1] ),
    .A(\top_inst.background_inst.counter_v[1] ),
    .X(_0280_));
 sg13g2_xnor2_1 _1871_ (.Y(_0281_),
    .A(_0479_),
    .B(_0280_));
 sg13g2_a21oi_2 _1872_ (.B1(_0281_),
    .Y(_0282_),
    .A2(_0279_),
    .A1(_0278_));
 sg13g2_xnor2_1 _1873_ (.Y(_0283_),
    .A(_0478_),
    .B(_0499_));
 sg13g2_xnor2_1 _1874_ (.Y(_0284_),
    .A(net42),
    .B(_0283_));
 sg13g2_a21oi_1 _1875_ (.A1(_0497_),
    .A2(_0555_),
    .Y(_0285_),
    .B1(_0479_));
 sg13g2_nor2_1 _1876_ (.A(_0228_),
    .B(_0285_),
    .Y(_0286_));
 sg13g2_a21o_1 _1877_ (.A2(_0284_),
    .A1(_0282_),
    .B1(_0286_),
    .X(_0287_));
 sg13g2_or2_1 _1878_ (.X(_0288_),
    .B(_0284_),
    .A(_0282_));
 sg13g2_nand4_1 _1879_ (.B(_0277_),
    .C(_0287_),
    .A(_0267_),
    .Y(_0289_),
    .D(_0288_));
 sg13g2_a21oi_1 _1880_ (.A1(_0271_),
    .A2(_0272_),
    .Y(_0290_),
    .B1(_0589_));
 sg13g2_o21ai_1 _1881_ (.B1(net36),
    .Y(_0291_),
    .A1(_0268_),
    .A2(_0290_));
 sg13g2_nand3_1 _1882_ (.B(_0271_),
    .C(_0272_),
    .A(_0589_),
    .Y(_0292_));
 sg13g2_nand2_1 _1883_ (.Y(_0293_),
    .A(_0268_),
    .B(_0292_));
 sg13g2_nand2_1 _1884_ (.Y(_0294_),
    .A(_0291_),
    .B(_0293_));
 sg13g2_a221oi_1 _1885_ (.B2(_0265_),
    .C1(net29),
    .B1(_0254_),
    .A1(_0260_),
    .Y(_0295_),
    .A2(_0261_));
 sg13g2_nand4_1 _1886_ (.B(_0260_),
    .C(_0261_),
    .A(net29),
    .Y(_0296_),
    .D(_0254_));
 sg13g2_nand3_1 _1887_ (.B(_0255_),
    .C(_0296_),
    .A(_0257_),
    .Y(_0297_));
 sg13g2_nand2b_1 _1888_ (.Y(_0298_),
    .B(_0297_),
    .A_N(_0295_));
 sg13g2_a21oi_1 _1889_ (.A1(_0494_),
    .A2(_0292_),
    .Y(_0299_),
    .B1(_0290_));
 sg13g2_nor2b_1 _1890_ (.A(_0299_),
    .B_N(_0268_),
    .Y(_0300_));
 sg13g2_a221oi_1 _1891_ (.B2(_0298_),
    .C1(_0300_),
    .B1(_0277_),
    .A1(net50),
    .Y(_0301_),
    .A2(_0294_));
 sg13g2_xnor2_1 _1892_ (.Y(_0302_),
    .A(_0507_),
    .B(\top_inst.background_inst.cur_time[7] ));
 sg13g2_xnor2_1 _1893_ (.Y(_0303_),
    .A(_0483_),
    .B(_0302_));
 sg13g2_o21ai_1 _1894_ (.B1(net49),
    .Y(_0304_),
    .A1(net46),
    .A2(_0583_));
 sg13g2_o21ai_1 _1895_ (.B1(_0304_),
    .Y(_0305_),
    .A1(_0722_),
    .A2(_0584_));
 sg13g2_xor2_1 _1896_ (.B(_0305_),
    .A(_0303_),
    .X(_0306_));
 sg13g2_nand2b_1 _1897_ (.Y(_0307_),
    .B(_0306_),
    .A_N(net44));
 sg13g2_a21oi_2 _1898_ (.B1(_0307_),
    .Y(_0308_),
    .A2(_0301_),
    .A1(_0289_));
 sg13g2_nor2_1 _1899_ (.A(\top_inst.background_inst.bg_select[0] ),
    .B(_0306_),
    .Y(_0309_));
 sg13g2_and3_1 _1900_ (.X(_0310_),
    .A(_0289_),
    .B(_0301_),
    .C(_0309_));
 sg13g2_buf_2 _1901_ (.A(_0310_),
    .X(_0311_));
 sg13g2_nor3_2 _1902_ (.A(_0250_),
    .B(_0308_),
    .C(_0311_),
    .Y(_0312_));
 sg13g2_xnor2_1 _1903_ (.Y(_0313_),
    .A(_0197_),
    .B(_0274_));
 sg13g2_xor2_1 _1904_ (.B(_0286_),
    .A(_0284_),
    .X(_0314_));
 sg13g2_nand3_1 _1905_ (.B(_0282_),
    .C(_0314_),
    .A(_0267_),
    .Y(_0315_));
 sg13g2_and3_1 _1906_ (.X(_0316_),
    .A(_0275_),
    .B(_0282_),
    .C(_0314_));
 sg13g2_a21oi_1 _1907_ (.A1(_0267_),
    .A2(_0316_),
    .Y(_0317_),
    .B1(_0273_));
 sg13g2_a21o_1 _1908_ (.A2(_0315_),
    .A1(_0313_),
    .B1(_0317_),
    .X(_0318_));
 sg13g2_nor3_1 _1909_ (.A(_0525_),
    .B(net41),
    .C(_0263_),
    .Y(_0319_));
 sg13g2_nor3_1 _1910_ (.A(_0525_),
    .B(net29),
    .C(_0259_),
    .Y(_0320_));
 sg13g2_o21ai_1 _1911_ (.B1(_0566_),
    .Y(_0321_),
    .A1(_0228_),
    .A2(_0285_));
 sg13g2_o21ai_1 _1912_ (.B1(_0321_),
    .Y(_0322_),
    .A1(_0319_),
    .A2(_0320_));
 sg13g2_nor3_1 _1913_ (.A(_0566_),
    .B(_0228_),
    .C(_0285_),
    .Y(_0323_));
 sg13g2_nor2_1 _1914_ (.A(_0525_),
    .B(_0233_),
    .Y(_0324_));
 sg13g2_nand2_1 _1915_ (.Y(_0325_),
    .A(_0478_),
    .B(net31));
 sg13g2_nor2_1 _1916_ (.A(\top_inst.background_inst.cur_time[3] ),
    .B(_0325_),
    .Y(_0326_));
 sg13g2_nor3_1 _1917_ (.A(net29),
    .B(_0259_),
    .C(_0325_),
    .Y(_0327_));
 sg13g2_a221oi_1 _1918_ (.B2(_0259_),
    .C1(_0327_),
    .B1(_0326_),
    .A1(_0323_),
    .Y(_0328_),
    .A2(_0324_));
 sg13g2_nand2_1 _1919_ (.Y(_0329_),
    .A(_0528_),
    .B(_0241_));
 sg13g2_nand2_1 _1920_ (.Y(_0330_),
    .A(_0496_),
    .B(net41));
 sg13g2_a22oi_1 _1921_ (.Y(_0331_),
    .B1(_0329_),
    .B2(_0330_),
    .A2(_0328_),
    .A1(_0322_));
 sg13g2_nand3_1 _1922_ (.B(_0496_),
    .C(net41),
    .A(_0528_),
    .Y(_0332_));
 sg13g2_xnor2_1 _1923_ (.Y(_0333_),
    .A(net41),
    .B(_0263_));
 sg13g2_nand2_1 _1924_ (.Y(_0334_),
    .A(_0257_),
    .B(_0333_));
 sg13g2_a21oi_1 _1925_ (.A1(_0735_),
    .A2(_0321_),
    .Y(_0335_),
    .B1(_0323_));
 sg13g2_a21oi_1 _1926_ (.A1(_0332_),
    .A2(_0334_),
    .Y(_0336_),
    .B1(_0335_));
 sg13g2_a21oi_1 _1927_ (.A1(_0330_),
    .A2(_0329_),
    .Y(_0337_),
    .B1(_0265_));
 sg13g2_a21oi_1 _1928_ (.A1(_0322_),
    .A2(_0328_),
    .Y(_0338_),
    .B1(_0265_));
 sg13g2_nor4_1 _1929_ (.A(_0331_),
    .B(_0336_),
    .C(_0337_),
    .D(_0338_),
    .Y(_0339_));
 sg13g2_nor2_1 _1930_ (.A(_0548_),
    .B(_0270_),
    .Y(_0340_));
 sg13g2_and2_1 _1931_ (.A(_0339_),
    .B(_0340_),
    .X(_0341_));
 sg13g2_nor4_1 _1932_ (.A(_0548_),
    .B(_0270_),
    .C(_0273_),
    .D(_0275_),
    .Y(_0342_));
 sg13g2_a21oi_2 _1933_ (.B1(_0342_),
    .Y(_0343_),
    .A2(_0341_),
    .A1(_0318_));
 sg13g2_a21oi_1 _1934_ (.A1(_0313_),
    .A2(_0315_),
    .Y(_0344_),
    .B1(_0317_));
 sg13g2_xor2_1 _1935_ (.B(_0269_),
    .A(_0268_),
    .X(_0345_));
 sg13g2_nor2_1 _1936_ (.A(net44),
    .B(_0345_),
    .Y(_0346_));
 sg13g2_nor2_1 _1937_ (.A(_0273_),
    .B(_0275_),
    .Y(_0347_));
 sg13g2_or3_1 _1938_ (.A(net44),
    .B(_0345_),
    .C(_0347_),
    .X(_0348_));
 sg13g2_nor2_1 _1939_ (.A(_0244_),
    .B(_0274_),
    .Y(_0349_));
 sg13g2_nand3_1 _1940_ (.B(_0241_),
    .C(_0349_),
    .A(_0239_),
    .Y(_0350_));
 sg13g2_o21ai_1 _1941_ (.B1(net44),
    .Y(_0351_),
    .A1(_0274_),
    .A2(_0271_));
 sg13g2_inv_1 _1942_ (.Y(_0352_),
    .A(_0351_));
 sg13g2_nand3_1 _1943_ (.B(net43),
    .C(_0552_),
    .A(net32),
    .Y(_0353_));
 sg13g2_a21oi_1 _1944_ (.A1(_0734_),
    .A2(_0552_),
    .Y(_0354_),
    .B1(net43));
 sg13g2_a221oi_1 _1945_ (.B2(_0897_),
    .C1(_0354_),
    .B1(_0353_),
    .A1(net29),
    .Y(_0355_),
    .A2(_0566_));
 sg13g2_nor3_1 _1946_ (.A(net31),
    .B(_0238_),
    .C(_0355_),
    .Y(_0356_));
 sg13g2_a21oi_1 _1947_ (.A1(_0897_),
    .A2(_0353_),
    .Y(_0357_),
    .B1(_0354_));
 sg13g2_nor3_1 _1948_ (.A(net42),
    .B(_0238_),
    .C(_0357_),
    .Y(_0358_));
 sg13g2_and2_1 _1949_ (.A(_0274_),
    .B(_0271_),
    .X(_0359_));
 sg13g2_o21ai_1 _1950_ (.B1(_0359_),
    .Y(_0360_),
    .A1(_0356_),
    .A2(_0358_));
 sg13g2_o21ai_1 _1951_ (.B1(_0206_),
    .Y(_0361_),
    .A1(net29),
    .A2(_0235_));
 sg13g2_a21oi_1 _1952_ (.A1(net33),
    .A2(_0361_),
    .Y(_0362_),
    .B1(_0889_));
 sg13g2_nor2_1 _1953_ (.A(net33),
    .B(_0361_),
    .Y(_0363_));
 sg13g2_o21ai_1 _1954_ (.B1(_0274_),
    .Y(_0364_),
    .A1(_0362_),
    .A2(_0363_));
 sg13g2_nand4_1 _1955_ (.B(_0352_),
    .C(_0360_),
    .A(_0350_),
    .Y(_0365_),
    .D(_0364_));
 sg13g2_o21ai_1 _1956_ (.B1(_0365_),
    .Y(_0366_),
    .A1(_0339_),
    .A2(_0348_));
 sg13g2_a21oi_2 _1957_ (.B1(_0366_),
    .Y(_0367_),
    .A2(_0346_),
    .A1(_0344_));
 sg13g2_nand2_2 _1958_ (.Y(_0368_),
    .A(_0343_),
    .B(_0367_));
 sg13g2_mux4_1 _1959_ (.S0(_0312_),
    .A0(_0221_),
    .A1(_0222_),
    .A2(_0223_),
    .A3(_0224_),
    .S1(_0368_),
    .X(_0369_));
 sg13g2_nor2_2 _1960_ (.A(\top_inst.background_inst.bg_select[1] ),
    .B(_0219_),
    .Y(_0370_));
 sg13g2_o21ai_1 _1961_ (.B1(_0240_),
    .Y(_0371_),
    .A1(_0566_),
    .A2(_0283_));
 sg13g2_xnor2_1 _1962_ (.Y(_0372_),
    .A(net50),
    .B(_0494_));
 sg13g2_nand2_1 _1963_ (.Y(_0373_),
    .A(_0372_),
    .B(_0256_));
 sg13g2_nand2_1 _1964_ (.Y(_0374_),
    .A(_0589_),
    .B(_0256_));
 sg13g2_nor3_1 _1965_ (.A(_0240_),
    .B(_0566_),
    .C(_0283_),
    .Y(_0375_));
 sg13g2_a221oi_1 _1966_ (.B2(_0374_),
    .C1(_0375_),
    .B1(_0373_),
    .A1(_0259_),
    .Y(_0376_),
    .A2(_0371_));
 sg13g2_nand2b_1 _1967_ (.Y(_0377_),
    .B(_0372_),
    .A_N(_0572_));
 sg13g2_a221oi_1 _1968_ (.B2(_0831_),
    .C1(_0375_),
    .B1(_0377_),
    .A1(_0259_),
    .Y(_0378_),
    .A2(_0371_));
 sg13g2_a22oi_1 _1969_ (.Y(_0379_),
    .B1(_0256_),
    .B2(_0585_),
    .A2(_0372_),
    .A1(_0589_));
 sg13g2_o21ai_1 _1970_ (.B1(_0379_),
    .Y(_0380_),
    .A1(_0572_),
    .A2(_0373_));
 sg13g2_nor3_2 _1971_ (.A(_0376_),
    .B(_0378_),
    .C(_0380_),
    .Y(_0381_));
 sg13g2_xor2_1 _1972_ (.B(net46),
    .A(net49),
    .X(_0382_));
 sg13g2_a21o_1 _1973_ (.A2(_0381_),
    .A1(_0583_),
    .B1(_0382_),
    .X(_0383_));
 sg13g2_o21ai_1 _1974_ (.B1(_0383_),
    .Y(_0384_),
    .A1(_0583_),
    .A2(_0381_));
 sg13g2_xor2_1 _1975_ (.B(_0384_),
    .A(_0303_),
    .X(_0385_));
 sg13g2_nor2_1 _1976_ (.A(net34),
    .B(\top_inst.background_inst.color3[5] ),
    .Y(_0386_));
 sg13g2_a21oi_1 _1977_ (.A1(net34),
    .A2(_0385_),
    .Y(_0387_),
    .B1(_0386_));
 sg13g2_nor2b_2 _1978_ (.A(_0731_),
    .B_N(_0218_),
    .Y(_0388_));
 sg13g2_nand3_1 _1979_ (.B(\top_inst.background_inst.color2[5] ),
    .C(net26),
    .A(_0212_),
    .Y(_0389_));
 sg13g2_o21ai_1 _1980_ (.B1(_0389_),
    .Y(_0390_),
    .A1(_0221_),
    .A2(net26));
 sg13g2_a22oi_1 _1981_ (.Y(_0391_),
    .B1(_0388_),
    .B2(_0390_),
    .A2(_0387_),
    .A1(_0370_));
 sg13g2_o21ai_1 _1982_ (.B1(_0391_),
    .Y(net8),
    .A1(_0220_),
    .A2(_0369_));
 sg13g2_nor2_1 _1983_ (.A(_0211_),
    .B(_0219_),
    .Y(_0392_));
 sg13g2_mux2_1 _1984_ (.A0(\top_inst.background_inst.color1[3] ),
    .A1(\top_inst.background_inst.color3[3] ),
    .S(_0312_),
    .X(_0393_));
 sg13g2_mux2_1 _1985_ (.A0(\top_inst.background_inst.color2[3] ),
    .A1(\top_inst.background_inst.color4[3] ),
    .S(_0312_),
    .X(_0394_));
 sg13g2_mux2_1 _1986_ (.A0(_0393_),
    .A1(_0394_),
    .S(_0368_),
    .X(_0395_));
 sg13g2_inv_1 _1987_ (.Y(_0396_),
    .A(\top_inst.background_inst.color1[3] ));
 sg13g2_nand3_1 _1988_ (.B(\top_inst.background_inst.color2[3] ),
    .C(_0738_),
    .A(_0212_),
    .Y(_0397_));
 sg13g2_o21ai_1 _1989_ (.B1(_0397_),
    .Y(_0398_),
    .A1(_0396_),
    .A2(_0739_));
 sg13g2_a21o_1 _1990_ (.A2(_0371_),
    .A1(_0259_),
    .B1(_0375_),
    .X(_0399_));
 sg13g2_inv_1 _1991_ (.Y(_0400_),
    .A(_0256_));
 sg13g2_a21o_1 _1992_ (.A2(_0399_),
    .A1(net33),
    .B1(_0400_),
    .X(_0401_));
 sg13g2_o21ai_1 _1993_ (.B1(_0401_),
    .Y(_0402_),
    .A1(net33),
    .A2(_0399_));
 sg13g2_xnor2_1 _1994_ (.Y(_0403_),
    .A(_0402_),
    .B(_0275_));
 sg13g2_nor2b_1 _1995_ (.A(net44),
    .B_N(\top_inst.background_inst.color3[3] ),
    .Y(_0404_));
 sg13g2_a21oi_1 _1996_ (.A1(net34),
    .A2(_0403_),
    .Y(_0405_),
    .B1(_0404_));
 sg13g2_nor3_1 _1997_ (.A(\top_inst.background_inst.bg_select[1] ),
    .B(_0219_),
    .C(_0405_),
    .Y(_0406_));
 sg13g2_a21o_1 _1998_ (.A2(_0398_),
    .A1(_0388_),
    .B1(_0406_),
    .X(_0407_));
 sg13g2_a21o_1 _1999_ (.A2(_0395_),
    .A1(_0392_),
    .B1(_0407_),
    .X(net9));
 sg13g2_inv_1 _2000_ (.Y(_0408_),
    .A(\top_inst.background_inst.color1[1] ));
 sg13g2_inv_1 _2001_ (.Y(_0409_),
    .A(\top_inst.background_inst.color3[1] ));
 sg13g2_inv_1 _2002_ (.Y(_0410_),
    .A(\top_inst.background_inst.color2[1] ));
 sg13g2_inv_1 _2003_ (.Y(_0411_),
    .A(\top_inst.background_inst.color4[1] ));
 sg13g2_mux4_1 _2004_ (.S0(_0312_),
    .A0(_0408_),
    .A1(_0409_),
    .A2(_0410_),
    .A3(_0411_),
    .S1(_0368_),
    .X(_0412_));
 sg13g2_nand3_1 _2005_ (.B(\top_inst.background_inst.color2[1] ),
    .C(_0738_),
    .A(_0212_),
    .Y(_0413_));
 sg13g2_o21ai_1 _2006_ (.B1(_0413_),
    .Y(_0414_),
    .A1(_0408_),
    .A2(net26));
 sg13g2_nor2_1 _2007_ (.A(_0566_),
    .B(_0283_),
    .Y(_0415_));
 sg13g2_xnor2_1 _2008_ (.Y(_0416_),
    .A(_0415_),
    .B(_0333_));
 sg13g2_nor2_1 _2009_ (.A(net34),
    .B(\top_inst.background_inst.color3[1] ),
    .Y(_0417_));
 sg13g2_a21oi_1 _2010_ (.A1(net34),
    .A2(_0416_),
    .Y(_0418_),
    .B1(_0417_));
 sg13g2_a22oi_1 _2011_ (.Y(_0419_),
    .B1(_0418_),
    .B2(_0370_),
    .A2(_0414_),
    .A1(_0388_));
 sg13g2_o21ai_1 _2012_ (.B1(_0419_),
    .Y(net10),
    .A1(_0220_),
    .A2(_0412_));
 sg13g2_nor4_1 _2013_ (.A(\top_inst.background_inst.color3[4] ),
    .B(_0250_),
    .C(_0308_),
    .D(_0311_),
    .Y(_0420_));
 sg13g2_nand3_1 _2014_ (.B(_0367_),
    .C(_0420_),
    .A(_0343_),
    .Y(_0421_));
 sg13g2_a21o_1 _2015_ (.A2(_0341_),
    .A1(_0318_),
    .B1(_0342_),
    .X(_0422_));
 sg13g2_buf_1 _2016_ (.A(_0422_),
    .X(_0423_));
 sg13g2_a21o_1 _2017_ (.A2(_0346_),
    .A1(_0344_),
    .B1(_0366_),
    .X(_0424_));
 sg13g2_buf_1 _2018_ (.A(_0424_),
    .X(_0425_));
 sg13g2_nor4_1 _2019_ (.A(\top_inst.background_inst.color4[4] ),
    .B(_0250_),
    .C(_0308_),
    .D(_0311_),
    .Y(_0426_));
 sg13g2_o21ai_1 _2020_ (.B1(_0426_),
    .Y(_0427_),
    .A1(_0423_),
    .A2(_0425_));
 sg13g2_nand3_1 _2021_ (.B(_0421_),
    .C(_0427_),
    .A(_0392_),
    .Y(_0428_));
 sg13g2_or3_1 _2022_ (.A(_0250_),
    .B(_0308_),
    .C(_0311_),
    .X(_0429_));
 sg13g2_o21ai_1 _2023_ (.B1(\top_inst.background_inst.color2[4] ),
    .Y(_0430_),
    .A1(_0423_),
    .A2(_0425_));
 sg13g2_nand3_1 _2024_ (.B(_0343_),
    .C(_0367_),
    .A(\top_inst.background_inst.color1[4] ),
    .Y(_0431_));
 sg13g2_and3_1 _2025_ (.X(_0432_),
    .A(_0429_),
    .B(_0430_),
    .C(_0431_));
 sg13g2_xnor2_1 _2026_ (.Y(_0433_),
    .A(_0381_),
    .B(_0268_));
 sg13g2_nor2_1 _2027_ (.A(net34),
    .B(\top_inst.background_inst.color3[4] ),
    .Y(_0434_));
 sg13g2_a21oi_1 _2028_ (.A1(_0549_),
    .A2(_0433_),
    .Y(_0435_),
    .B1(_0434_));
 sg13g2_inv_1 _2029_ (.Y(_0436_),
    .A(\top_inst.background_inst.color1[4] ));
 sg13g2_nand3_1 _2030_ (.B(\top_inst.background_inst.color2[4] ),
    .C(net26),
    .A(_0212_),
    .Y(_0437_));
 sg13g2_o21ai_1 _2031_ (.B1(_0437_),
    .Y(_0438_),
    .A1(_0436_),
    .A2(net26));
 sg13g2_a22oi_1 _2032_ (.Y(_0439_),
    .B1(_0438_),
    .B2(_0388_),
    .A2(_0435_),
    .A1(_0370_));
 sg13g2_o21ai_1 _2033_ (.B1(_0439_),
    .Y(net12),
    .A1(_0428_),
    .A2(_0432_));
 sg13g2_nor4_1 _2034_ (.A(\top_inst.background_inst.color3[2] ),
    .B(_0250_),
    .C(_0308_),
    .D(_0311_),
    .Y(_0440_));
 sg13g2_nand3_1 _2035_ (.B(_0367_),
    .C(_0440_),
    .A(_0343_),
    .Y(_0441_));
 sg13g2_nor4_1 _2036_ (.A(\top_inst.background_inst.color4[2] ),
    .B(_0250_),
    .C(_0308_),
    .D(_0311_),
    .Y(_0442_));
 sg13g2_o21ai_1 _2037_ (.B1(_0442_),
    .Y(_0443_),
    .A1(_0423_),
    .A2(_0425_));
 sg13g2_nand3_1 _2038_ (.B(_0441_),
    .C(_0443_),
    .A(_0392_),
    .Y(_0444_));
 sg13g2_o21ai_1 _2039_ (.B1(\top_inst.background_inst.color2[2] ),
    .Y(_0445_),
    .A1(_0423_),
    .A2(_0425_));
 sg13g2_nand3_1 _2040_ (.B(_0343_),
    .C(_0367_),
    .A(\top_inst.background_inst.color1[2] ),
    .Y(_0446_));
 sg13g2_and3_1 _2041_ (.X(_0447_),
    .A(_0429_),
    .B(_0445_),
    .C(_0446_));
 sg13g2_xnor2_1 _2042_ (.Y(_0448_),
    .A(_0399_),
    .B(_0257_));
 sg13g2_nor2_1 _2043_ (.A(net34),
    .B(\top_inst.background_inst.color3[2] ),
    .Y(_0449_));
 sg13g2_a21oi_1 _2044_ (.A1(_0549_),
    .A2(_0448_),
    .Y(_0450_),
    .B1(_0449_));
 sg13g2_inv_1 _2045_ (.Y(_0451_),
    .A(\top_inst.background_inst.color1[2] ));
 sg13g2_nand3_1 _2046_ (.B(\top_inst.background_inst.color2[2] ),
    .C(net26),
    .A(_0212_),
    .Y(_0452_));
 sg13g2_o21ai_1 _2047_ (.B1(_0452_),
    .Y(_0453_),
    .A1(_0451_),
    .A2(net26));
 sg13g2_a22oi_1 _2048_ (.Y(_0454_),
    .B1(_0453_),
    .B2(_0388_),
    .A2(_0450_),
    .A1(_0370_));
 sg13g2_o21ai_1 _2049_ (.B1(_0454_),
    .Y(net13),
    .A1(_0444_),
    .A2(_0447_));
 sg13g2_nor2b_1 _2050_ (.A(net44),
    .B_N(\top_inst.background_inst.color3[0] ),
    .Y(_0455_));
 sg13g2_a21oi_1 _2051_ (.A1(net44),
    .A2(_0284_),
    .Y(_0456_),
    .B1(_0455_));
 sg13g2_nor2_1 _2052_ (.A(\top_inst.background_inst.bg_select[1] ),
    .B(_0456_),
    .Y(_0457_));
 sg13g2_or3_1 _2053_ (.A(\top_inst.background_inst.color1[0] ),
    .B(_0312_),
    .C(_0457_),
    .X(_0458_));
 sg13g2_nand2_1 _2054_ (.Y(_0459_),
    .A(_0212_),
    .B(_0738_));
 sg13g2_nand2b_1 _2055_ (.Y(_0460_),
    .B(_0737_),
    .A_N(\top_inst.background_inst.color1[0] ));
 sg13g2_a21oi_1 _2056_ (.A1(_0459_),
    .A2(_0460_),
    .Y(_0461_),
    .B1(_0731_));
 sg13g2_nor2b_1 _2057_ (.A(_0461_),
    .B_N(_0218_),
    .Y(_0462_));
 sg13g2_o21ai_1 _2058_ (.B1(_0462_),
    .Y(_0463_),
    .A1(_0368_),
    .A2(_0458_));
 sg13g2_nand2b_1 _2059_ (.Y(_0464_),
    .B(_0312_),
    .A_N(\top_inst.background_inst.color3[0] ));
 sg13g2_nor3_1 _2060_ (.A(_0211_),
    .B(_0423_),
    .C(_0425_),
    .Y(_0465_));
 sg13g2_a21oi_1 _2061_ (.A1(_0343_),
    .A2(_0367_),
    .Y(_0466_),
    .B1(_0211_));
 sg13g2_mux2_1 _2062_ (.A0(\top_inst.background_inst.color4[0] ),
    .A1(\top_inst.background_inst.color2[0] ),
    .S(_0429_),
    .X(_0467_));
 sg13g2_nor2_1 _2063_ (.A(_0731_),
    .B(_0738_),
    .Y(_0468_));
 sg13g2_or2_1 _2064_ (.X(_0469_),
    .B(_0468_),
    .A(_0457_));
 sg13g2_a221oi_1 _2065_ (.B2(_0467_),
    .C1(_0469_),
    .B1(_0466_),
    .A1(_0464_),
    .Y(_0470_),
    .A2(_0465_));
 sg13g2_nand4_1 _2066_ (.B(_0212_),
    .C(net26),
    .A(\top_inst.background_inst.color2[0] ),
    .Y(_0471_),
    .D(_0388_));
 sg13g2_o21ai_1 _2067_ (.B1(_0471_),
    .Y(net14),
    .A1(_0463_),
    .A2(_0470_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _2072__107 (.L_HI(net107));
 sg13g2_buf_1 _2070_ (.A(net96),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2071_ (.A(net97),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2072_ (.A(net107),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2073_ (.A(net98),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2074_ (.A(net108),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2075_ (.A(net109),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2076_ (.A(net99),
    .X(uio_oe[6]));
 sg13g2_buf_1 _2077_ (.A(net100),
    .X(uio_oe[7]));
 sg13g2_buf_1 _2078_ (.A(net101),
    .X(uio_out[0]));
 sg13g2_buf_1 _2079_ (.A(net102),
    .X(uio_out[1]));
 sg13g2_buf_1 _2080_ (.A(net103),
    .X(uio_out[2]));
 sg13g2_buf_1 _2081_ (.A(net104),
    .X(uio_out[3]));
 sg13g2_buf_1 _2082_ (.A(net23),
    .X(net6));
 sg13g2_buf_1 _2083_ (.A(net19),
    .X(net7));
 sg13g2_buf_1 _2084_ (.A(net105),
    .X(uio_out[6]));
 sg13g2_buf_1 _2085_ (.A(net106),
    .X(uio_out[7]));
 sg13g2_buf_1 _2086_ (.A(\top_inst.timing_ver.sync ),
    .X(net11));
 sg13g2_buf_1 _2087_ (.A(hsync),
    .X(net15));
 sg13g2_dfrbp_1 \top_inst.bg_sel[0]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_1351_clk),
    .RESET_B(net91),
    .D(_0102_),
    .Q_N(_1017_),
    .Q(\top_inst.background_inst.bg_select[0] ));
 sg13g2_dfrbp_1 \top_inst.bg_sel[1]$_DFFE_PN1P_  (.CLK(clknet_level_3_1_1351_clk),
    .RESET_B(net73),
    .D(_0103_),
    .Q_N(\top_inst.background_inst.bg_select[1] ),
    .Q(_0047_));
 sg13g2_dfrbp_1 \top_inst.cur_time[0]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_1247_clk),
    .RESET_B(net92),
    .D(_0104_),
    .Q_N(_0043_),
    .Q(\top_inst.background_inst.cur_time[0] ));
 sg13g2_dfrbp_1 \top_inst.cur_time[1]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_1247_clk),
    .RESET_B(net92),
    .D(_0105_),
    .Q_N(_1016_),
    .Q(\top_inst.background_inst.cur_time[1] ));
 sg13g2_dfrbp_1 \top_inst.cur_time[2]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_1559_clk),
    .RESET_B(net92),
    .D(_0106_),
    .Q_N(_1015_),
    .Q(\top_inst.background_inst.cur_time[2] ));
 sg13g2_dfrbp_1 \top_inst.cur_time[3]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_1559_clk),
    .RESET_B(net92),
    .D(_0107_),
    .Q_N(_1014_),
    .Q(\top_inst.background_inst.cur_time[3] ));
 sg13g2_dfrbp_1 \top_inst.cur_time[4]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_1455_clk),
    .RESET_B(net93),
    .D(_0108_),
    .Q_N(_1013_),
    .Q(\top_inst.background_inst.cur_time[4] ));
 sg13g2_dfrbp_1 \top_inst.cur_time[5]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_1559_clk),
    .RESET_B(net93),
    .D(_0109_),
    .Q_N(_1012_),
    .Q(\top_inst.background_inst.cur_time[5] ));
 sg13g2_dfrbp_1 \top_inst.cur_time[6]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_1247_clk),
    .RESET_B(net92),
    .D(_0110_),
    .Q_N(_1011_),
    .Q(\top_inst.background_inst.cur_time[6] ));
 sg13g2_dfrbp_1 \top_inst.cur_time[7]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_1247_clk),
    .RESET_B(net92),
    .D(_0111_),
    .Q_N(_1018_),
    .Q(\top_inst.background_inst.cur_time[7] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.load_register$_DFF_PN0_  (.CLK(clknet_level_3_1_623_clk),
    .RESET_B(net68),
    .D(_0012_),
    .Q_N(_1010_),
    .Q(\top_inst.spi_receiver_inst.load_register ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[0][0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0000_),
    .GATE_N(clknet_1_0__leaf__0021_),
    .RESET_B(net110),
    .Q(\top_inst.background_inst.color1[0] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[0][1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0001_),
    .GATE_N(clknet_1_1__leaf__0021_),
    .RESET_B(net111),
    .Q(\top_inst.background_inst.color1[1] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[0][2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0002_),
    .GATE_N(clknet_1_0__leaf__0021_),
    .RESET_B(net112),
    .Q(\top_inst.background_inst.color1[2] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[0][3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0003_),
    .GATE_N(clknet_1_1__leaf__0021_),
    .RESET_B(net113),
    .Q(\top_inst.background_inst.color1[3] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[0][4]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0004_),
    .GATE_N(clknet_1_1__leaf__0021_),
    .RESET_B(net114),
    .Q(\top_inst.background_inst.color1[4] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[0][5]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0005_),
    .GATE_N(clknet_1_0__leaf__0021_),
    .RESET_B(net115),
    .Q(\top_inst.background_inst.color1[5] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[1][0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0000_),
    .GATE_N(clknet_1_0__leaf__0020_),
    .RESET_B(net116),
    .Q(\top_inst.background_inst.color2[0] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[1][1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0001_),
    .GATE_N(clknet_1_1__leaf__0020_),
    .RESET_B(net117),
    .Q(\top_inst.background_inst.color2[1] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[1][2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0006_),
    .GATE_N(clknet_1_1__leaf__0020_),
    .RESET_B(net118),
    .Q(\top_inst.background_inst.color2[2] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[1][3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0003_),
    .GATE_N(clknet_1_1__leaf__0020_),
    .RESET_B(net119),
    .Q(\top_inst.background_inst.color2[3] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[1][4]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0004_),
    .GATE_N(clknet_1_0__leaf__0020_),
    .RESET_B(net120),
    .Q(\top_inst.background_inst.color2[4] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[1][5]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0007_),
    .GATE_N(clknet_1_0__leaf__0020_),
    .RESET_B(net121),
    .Q(\top_inst.background_inst.color2[5] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[2][0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0008_),
    .GATE_N(clknet_1_0__leaf__0019_),
    .RESET_B(net122),
    .Q(\top_inst.background_inst.color3[0] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[2][1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0001_),
    .GATE_N(clknet_1_1__leaf__0019_),
    .RESET_B(net123),
    .Q(\top_inst.background_inst.color3[1] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[2][2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0006_),
    .GATE_N(clknet_1_0__leaf__0019_),
    .RESET_B(net124),
    .Q(\top_inst.background_inst.color3[2] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[2][3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0009_),
    .GATE_N(clknet_1_1__leaf__0019_),
    .RESET_B(net125),
    .Q(\top_inst.background_inst.color3[3] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[2][4]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0010_),
    .GATE_N(clknet_1_0__leaf__0019_),
    .RESET_B(net126),
    .Q(\top_inst.background_inst.color3[4] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[2][5]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0007_),
    .GATE_N(clknet_1_1__leaf__0019_),
    .RESET_B(net127),
    .Q(\top_inst.background_inst.color3[5] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[3][0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0008_),
    .GATE_N(clknet_1_0__leaf__0018_),
    .RESET_B(net128),
    .Q(\top_inst.background_inst.color4[0] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[3][1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0001_),
    .GATE_N(clknet_1_1__leaf__0018_),
    .RESET_B(net129),
    .Q(\top_inst.background_inst.color4[1] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[3][2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0006_),
    .GATE_N(clknet_1_1__leaf__0018_),
    .RESET_B(net130),
    .Q(\top_inst.background_inst.color4[2] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[3][3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0009_),
    .GATE_N(clknet_1_0__leaf__0018_),
    .RESET_B(net131),
    .Q(\top_inst.background_inst.color4[3] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[3][4]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0010_),
    .GATE_N(clknet_1_1__leaf__0018_),
    .RESET_B(net132),
    .Q(\top_inst.background_inst.color4[4] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[3][5]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0005_),
    .GATE_N(clknet_1_0__leaf__0018_),
    .RESET_B(net133),
    .Q(\top_inst.background_inst.color4[5] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[4][0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0008_),
    .GATE_N(clknet_1_0__leaf__0017_),
    .RESET_B(net134),
    .Q(\top_inst.spi_receiver_inst.registers[4][0] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[4][1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0001_),
    .GATE_N(clknet_1_1__leaf__0017_),
    .RESET_B(net135),
    .Q(\top_inst.spi_receiver_inst.registers[4][1] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[4][2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0002_),
    .GATE_N(clknet_1_1__leaf__0017_),
    .RESET_B(net136),
    .Q(\top_inst.spi_receiver_inst.registers[4][2] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[4][3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0003_),
    .GATE_N(clknet_1_1__leaf__0017_),
    .RESET_B(net137),
    .Q(\top_inst.spi_receiver_inst.registers[4][3] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[4][4]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0010_),
    .GATE_N(clknet_1_1__leaf__0017_),
    .RESET_B(net138),
    .Q(\top_inst.spi_receiver_inst.registers[4][4] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[4][5]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0007_),
    .GATE_N(clknet_1_0__leaf__0017_),
    .RESET_B(net139),
    .Q(\top_inst.spi_receiver_inst.registers[4][5] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[4][6]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0013_),
    .GATE_N(clknet_1_0__leaf__0017_),
    .RESET_B(net140),
    .Q(\top_inst.spi_receiver_inst.registers[4][6] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[4][7]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0014_),
    .GATE_N(clknet_1_0__leaf__0017_),
    .RESET_B(net141),
    .Q(\top_inst.spi_receiver_inst.registers[4][7] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[5][0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0008_),
    .GATE_N(clknet_1_0__leaf__0016_),
    .RESET_B(net142),
    .Q(\top_inst.spi_receiver_inst.registers[5][0] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[5][1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0001_),
    .GATE_N(clknet_1_1__leaf__0016_),
    .RESET_B(net143),
    .Q(\top_inst.spi_receiver_inst.registers[5][1] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[5][2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0002_),
    .GATE_N(clknet_1_1__leaf__0016_),
    .RESET_B(net144),
    .Q(\top_inst.spi_receiver_inst.registers[5][2] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[5][3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0003_),
    .GATE_N(clknet_1_1__leaf__0016_),
    .RESET_B(net145),
    .Q(\top_inst.spi_receiver_inst.registers[5][3] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[5][4]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0010_),
    .GATE_N(clknet_1_1__leaf__0016_),
    .RESET_B(net146),
    .Q(\top_inst.spi_receiver_inst.registers[5][4] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[5][5]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0007_),
    .GATE_N(clknet_1_0__leaf__0016_),
    .RESET_B(net147),
    .Q(\top_inst.spi_receiver_inst.registers[5][5] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[5][6]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0013_),
    .GATE_N(clknet_1_0__leaf__0016_),
    .RESET_B(net148),
    .Q(\top_inst.spi_receiver_inst.registers[5][6] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[5][7]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0014_),
    .GATE_N(clknet_1_0__leaf__0016_),
    .RESET_B(net149),
    .Q(\top_inst.spi_receiver_inst.registers[5][7] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[6][0]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0008_),
    .GATE_N(clknet_1_0__leaf__0015_),
    .RESET_B(net150),
    .Q(\top_inst.misc[0] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[6][1]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0011_),
    .GATE_N(clknet_1_0__leaf__0015_),
    .RESET_B(net151),
    .Q(\top_inst.misc[1] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[6][2]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0006_),
    .GATE_N(clknet_1_1__leaf__0015_),
    .RESET_B(net152),
    .Q(\top_inst.misc[2] ));
 sg13g2_dllrq_1 \top_inst.spi_receiver_inst.registers[6][3]$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(_0003_),
    .GATE_N(clknet_1_1__leaf__0015_),
    .RESET_B(net153),
    .Q(\top_inst.misc[3] ));
 sg13g2_lgcp_1 \top_inst.spi_receiver_inst.regs[0].sg13g2_lgcp_1_inst  (.GATE(_0022_),
    .CLK(clknet_level_3_1_831_clk),
    .GCLK(\top_inst.spi_receiver_inst.reg_gclk[0] ));
 sg13g2_lgcp_1 \top_inst.spi_receiver_inst.regs[1].sg13g2_lgcp_1_inst  (.GATE(_0023_),
    .CLK(clknet_level_3_1_727_clk),
    .GCLK(\top_inst.spi_receiver_inst.reg_gclk[1] ));
 sg13g2_lgcp_1 \top_inst.spi_receiver_inst.regs[2].sg13g2_lgcp_1_inst  (.GATE(_0024_),
    .CLK(clknet_level_3_1_727_clk),
    .GCLK(\top_inst.spi_receiver_inst.reg_gclk[2] ));
 sg13g2_lgcp_1 \top_inst.spi_receiver_inst.regs[3].sg13g2_lgcp_1_inst  (.GATE(_0025_),
    .CLK(clknet_level_3_1_727_clk),
    .GCLK(\top_inst.spi_receiver_inst.reg_gclk[3] ));
 sg13g2_lgcp_1 \top_inst.spi_receiver_inst.regs[4].sg13g2_lgcp_1_inst  (.GATE(_0026_),
    .CLK(clknet_level_3_1_623_clk),
    .GCLK(\top_inst.spi_receiver_inst.reg_gclk[4] ));
 sg13g2_lgcp_1 \top_inst.spi_receiver_inst.regs[5].sg13g2_lgcp_1_inst  (.GATE(_0027_),
    .CLK(clknet_level_3_1_623_clk),
    .GCLK(\top_inst.spi_receiver_inst.reg_gclk[5] ));
 sg13g2_lgcp_1 \top_inst.spi_receiver_inst.regs[6].sg13g2_lgcp_1_inst  (.GATE(_0028_),
    .CLK(clknet_level_3_1_727_clk),
    .GCLK(\top_inst.spi_receiver_inst.reg_gclk[6] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.spi_cmd[0]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_623_clk),
    .RESET_B(net70),
    .D(_0112_),
    .Q_N(_1009_),
    .Q(\top_inst.spi_receiver_inst.spi_cmd[0] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.spi_cmd[1]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_831_clk),
    .RESET_B(net68),
    .D(_0113_),
    .Q_N(_1008_),
    .Q(\top_inst.spi_receiver_inst.spi_cmd[1] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.spi_cmd[2]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_831_clk),
    .RESET_B(net68),
    .D(_0114_),
    .Q_N(_0041_),
    .Q(\top_inst.spi_receiver_inst.spi_cmd[2] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.spi_cnt[0]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_831_clk),
    .RESET_B(net69),
    .D(_0115_),
    .Q_N(_0044_),
    .Q(\top_inst.spi_receiver_inst.spi_cnt[0] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.spi_cnt[1]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_519_clk),
    .RESET_B(net68),
    .D(_0116_),
    .Q_N(_1007_),
    .Q(\top_inst.spi_receiver_inst.spi_cnt[1] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.spi_cnt[2]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_831_clk),
    .RESET_B(net69),
    .D(_0117_),
    .Q_N(_1006_),
    .Q(\top_inst.spi_receiver_inst.spi_cnt[2] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.spi_data[0]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_623_clk),
    .RESET_B(net69),
    .D(_0118_),
    .Q_N(_1005_),
    .Q(\top_inst.spi_receiver_inst.spi_data[0] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.spi_data[1]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_623_clk),
    .RESET_B(net70),
    .D(_0119_),
    .Q_N(_1004_),
    .Q(\top_inst.spi_receiver_inst.spi_data[1] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.spi_data[2]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_727_clk),
    .RESET_B(net73),
    .D(_0120_),
    .Q_N(_1003_),
    .Q(\top_inst.spi_receiver_inst.spi_data[2] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.spi_data[3]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_727_clk),
    .RESET_B(net73),
    .D(_0121_),
    .Q_N(_1002_),
    .Q(\top_inst.spi_receiver_inst.spi_data[3] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.spi_data[4]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_623_clk),
    .RESET_B(net70),
    .D(_0122_),
    .Q_N(_1001_),
    .Q(\top_inst.spi_receiver_inst.spi_data[4] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.spi_data[5]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_519_clk),
    .RESET_B(net69),
    .D(_0123_),
    .Q_N(_1000_),
    .Q(\top_inst.spi_receiver_inst.spi_data[5] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.spi_data[6]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_831_clk),
    .RESET_B(net68),
    .D(_0124_),
    .Q_N(_0999_),
    .Q(\top_inst.spi_receiver_inst.spi_data[6] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.spi_data[7]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_519_clk),
    .RESET_B(net68),
    .D(_0125_),
    .Q_N(_0998_),
    .Q(\top_inst.spi_receiver_inst.spi_data[7] ));
 sg13g2_dfrbp_1 \top_inst.spi_receiver_inst.spi_mode$_DFFE_PN0P_  (.CLK(clknet_level_3_1_831_clk),
    .RESET_B(net69),
    .D(_0126_),
    .Q_N(_1019_),
    .Q(\top_inst.spi_receiver_inst.spi_mode ));
 sg13g2_dfrbp_1 \top_inst.spi_sclk_delayed$_DFF_P_  (.CLK(clknet_level_3_1_1455_clk),
    .RESET_B(net154),
    .D(\top_inst.spi_receiver_inst.spi_sclk ),
    .Q_N(_0997_),
    .Q(\top_inst.spi_receiver_inst.spi_sclk_delayed ));
 sg13g2_dfrbp_1 \top_inst.sprite_access_inst.sprite_line[0]$_DFFE_PP_  (.CLK(clknet_level_3_1_1455_clk),
    .RESET_B(net155),
    .D(_0127_),
    .Q_N(_0996_),
    .Q(\top_inst.sprite_access_inst.sprite_line[0] ));
 sg13g2_dfrbp_1 \top_inst.sprite_access_inst.sprite_line[10]$_DFFE_PP_  (.CLK(clknet_level_3_1_1663_clk),
    .RESET_B(net156),
    .D(_0128_),
    .Q_N(_0995_),
    .Q(\top_inst.sprite_access_inst.sprite_line[10] ));
 sg13g2_dfrbp_1 \top_inst.sprite_access_inst.sprite_line[11]$_DFFE_PP_  (.CLK(clknet_level_3_1_1455_clk),
    .RESET_B(net157),
    .D(_0129_),
    .Q_N(_0994_),
    .Q(\top_inst.sprite_access_inst.sprite_line[11] ));
 sg13g2_dfrbp_1 \top_inst.sprite_access_inst.sprite_line[1]$_DFFE_PP_  (.CLK(clknet_level_3_1_1663_clk),
    .RESET_B(net158),
    .D(_0130_),
    .Q_N(_0993_),
    .Q(\top_inst.sprite_access_inst.sprite_line[1] ));
 sg13g2_dfrbp_1 \top_inst.sprite_access_inst.sprite_line[2]$_DFFE_PP_  (.CLK(clknet_level_3_1_1663_clk),
    .RESET_B(net159),
    .D(_0131_),
    .Q_N(_0992_),
    .Q(\top_inst.sprite_access_inst.sprite_line[2] ));
 sg13g2_dfrbp_1 \top_inst.sprite_access_inst.sprite_line[3]$_DFFE_PP_  (.CLK(clknet_level_3_1_1663_clk),
    .RESET_B(net160),
    .D(_0132_),
    .Q_N(_0991_),
    .Q(\top_inst.sprite_access_inst.sprite_line[3] ));
 sg13g2_dfrbp_1 \top_inst.sprite_access_inst.sprite_line[4]$_DFFE_PP_  (.CLK(clknet_level_3_1_1559_clk),
    .RESET_B(net161),
    .D(_0133_),
    .Q_N(_0990_),
    .Q(\top_inst.sprite_access_inst.sprite_line[4] ));
 sg13g2_dfrbp_1 \top_inst.sprite_access_inst.sprite_line[5]$_DFFE_PP_  (.CLK(clknet_level_3_1_1559_clk),
    .RESET_B(net162),
    .D(_0134_),
    .Q_N(_0989_),
    .Q(\top_inst.sprite_access_inst.sprite_line[5] ));
 sg13g2_dfrbp_1 \top_inst.sprite_access_inst.sprite_line[6]$_DFFE_PP_  (.CLK(clknet_level_3_1_1559_clk),
    .RESET_B(net163),
    .D(_0135_),
    .Q_N(_0988_),
    .Q(\top_inst.sprite_access_inst.sprite_line[6] ));
 sg13g2_dfrbp_1 \top_inst.sprite_access_inst.sprite_line[7]$_DFFE_PP_  (.CLK(clknet_level_3_1_1559_clk),
    .RESET_B(net164),
    .D(_0136_),
    .Q_N(_0987_),
    .Q(\top_inst.sprite_access_inst.sprite_line[7] ));
 sg13g2_dfrbp_1 \top_inst.sprite_access_inst.sprite_line[8]$_DFFE_PP_  (.CLK(clknet_level_3_1_1663_clk),
    .RESET_B(net165),
    .D(_0137_),
    .Q_N(_0986_),
    .Q(\top_inst.sprite_access_inst.sprite_line[8] ));
 sg13g2_dfrbp_1 \top_inst.sprite_access_inst.sprite_line[9]$_DFFE_PP_  (.CLK(clknet_level_3_1_1455_clk),
    .RESET_B(net166),
    .D(_0138_),
    .Q_N(_1020_),
    .Q(\top_inst.sprite_access_inst.sprite_line[9] ));
 sg13g2_lgcp_1 \top_inst.sprite_data_inst.sg13g2_lgcp_1_inst  (.GATE(\top_inst.sprite_data_inst.shiftf ),
    .CLK(clknet_4_10_0_clk),
    .GCLK(\top_inst.sprite_data_inst.gclk ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[0]$_DFF_PN0_  (.CLK(\clknet_5_31__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net89),
    .D(\top_inst.sprite_data_inst.sprite_data[1] ),
    .Q_N(_0985_),
    .Q(\top_inst.sprite_access_inst.sprite_data ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[100]$_DFF_PN1_  (.CLK(\clknet_5_23__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net85),
    .D(_0984_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[100] ),
    .Q(_1078_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[101]$_DFF_PN0_  (.CLK(\clknet_5_21__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net85),
    .D(\top_inst.sprite_data_inst.sprite_data[102] ),
    .Q_N(_0984_),
    .Q(\top_inst.sprite_data_inst.sprite_data[101] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[102]$_DFF_PN1_  (.CLK(\clknet_5_23__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net85),
    .D(_0055_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[102] ),
    .Q(_1079_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[103]$_DFF_PN1_  (.CLK(\clknet_5_21__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net85),
    .D(_1021_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[103] ),
    .Q(_1080_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[104]$_DFF_PN0_  (.CLK(\clknet_5_21__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net85),
    .D(\top_inst.sprite_data_inst.sprite_data[105] ),
    .Q_N(_1021_),
    .Q(\top_inst.sprite_data_inst.sprite_data[104] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[105]$_DFF_PN0_  (.CLK(\clknet_5_21__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net85),
    .D(\top_inst.sprite_data_inst.sprite_data[106] ),
    .Q_N(_1022_),
    .Q(\top_inst.sprite_data_inst.sprite_data[105] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[106]$_DFF_PN0_  (.CLK(\clknet_5_23__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net83),
    .D(\top_inst.sprite_data_inst.sprite_data[107] ),
    .Q_N(_0983_),
    .Q(\top_inst.sprite_data_inst.sprite_data[106] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[107]$_DFF_PN1_  (.CLK(\clknet_5_20__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net83),
    .D(_0982_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[107] ),
    .Q(_1081_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[108]$_DFF_PN0_  (.CLK(\clknet_5_20__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net83),
    .D(\top_inst.sprite_data_inst.sprite_data[109] ),
    .Q_N(_0982_),
    .Q(\top_inst.sprite_data_inst.sprite_data[108] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[109]$_DFF_PN1_  (.CLK(\clknet_5_20__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net83),
    .D(_1024_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[109] ),
    .Q(_1082_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[10]$_DFF_PN0_  (.CLK(\clknet_5_27__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net88),
    .D(\top_inst.sprite_data_inst.sprite_data[11] ),
    .Q_N(_1023_),
    .Q(\top_inst.sprite_data_inst.sprite_data[10] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[110]$_DFF_PN0_  (.CLK(\clknet_5_19__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net77),
    .D(\top_inst.sprite_data_inst.sprite_data[111] ),
    .Q_N(_1024_),
    .Q(\top_inst.sprite_data_inst.sprite_data[110] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[111]$_DFF_PN0_  (.CLK(\clknet_5_17__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net77),
    .D(\top_inst.sprite_data_inst.sprite_data[112] ),
    .Q_N(_1025_),
    .Q(\top_inst.sprite_data_inst.sprite_data[111] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[112]$_DFF_PN0_  (.CLK(\clknet_5_17__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net77),
    .D(\top_inst.sprite_data_inst.sprite_data[113] ),
    .Q_N(_1026_),
    .Q(\top_inst.sprite_data_inst.sprite_data[112] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[113]$_DFF_PN0_  (.CLK(\clknet_5_17__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net77),
    .D(\top_inst.sprite_data_inst.sprite_data[114] ),
    .Q_N(_0981_),
    .Q(\top_inst.sprite_data_inst.sprite_data[113] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[114]$_DFF_PN1_  (.CLK(\clknet_5_16__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net75),
    .D(_0056_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[114] ),
    .Q(_1083_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[115]$_DFF_PN1_  (.CLK(\clknet_5_16__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net75),
    .D(_1027_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[115] ),
    .Q(_1084_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[116]$_DFF_PN0_  (.CLK(\clknet_5_16__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net75),
    .D(\top_inst.sprite_data_inst.sprite_data[117] ),
    .Q_N(_1027_),
    .Q(\top_inst.sprite_data_inst.sprite_data[116] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[117]$_DFF_PN0_  (.CLK(\clknet_5_22__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net83),
    .D(\top_inst.sprite_data_inst.sprite_data[118] ),
    .Q_N(_0980_),
    .Q(\top_inst.sprite_data_inst.sprite_data[117] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[118]$_DFF_PN1_  (.CLK(\clknet_5_20__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net83),
    .D(_1028_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[118] ),
    .Q(_1085_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[119]$_DFF_PN0_  (.CLK(\clknet_5_19__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net83),
    .D(\top_inst.sprite_data_inst.sprite_data[120] ),
    .Q_N(_1028_),
    .Q(\top_inst.sprite_data_inst.sprite_data[119] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[11]$_DFF_PN0_  (.CLK(\clknet_5_26__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net88),
    .D(\top_inst.sprite_data_inst.sprite_data[12] ),
    .Q_N(_1029_),
    .Q(\top_inst.sprite_data_inst.sprite_data[11] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[120]$_DFF_PN0_  (.CLK(\clknet_5_19__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net77),
    .D(\top_inst.sprite_data_inst.sprite_data[121] ),
    .Q_N(_1030_),
    .Q(\top_inst.sprite_data_inst.sprite_data[120] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[121]$_DFF_PN0_  (.CLK(\clknet_5_18__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net78),
    .D(\top_inst.sprite_data_inst.sprite_data[122] ),
    .Q_N(_0979_),
    .Q(\top_inst.sprite_data_inst.sprite_data[121] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[122]$_DFF_PN1_  (.CLK(\clknet_5_16__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net77),
    .D(_1031_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[122] ),
    .Q(_1086_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[123]$_DFF_PN0_  (.CLK(\clknet_5_18__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net77),
    .D(\top_inst.sprite_data_inst.sprite_data[124] ),
    .Q_N(_1031_),
    .Q(\top_inst.sprite_data_inst.sprite_data[123] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[124]$_DFF_PN0_  (.CLK(\clknet_5_7__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net75),
    .D(\top_inst.sprite_data_inst.sprite_data[125] ),
    .Q_N(_1032_),
    .Q(\top_inst.sprite_data_inst.sprite_data[124] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[125]$_DFF_PN0_  (.CLK(\clknet_5_7__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net76),
    .D(\top_inst.sprite_data_inst.sprite_data[126] ),
    .Q_N(_0978_),
    .Q(\top_inst.sprite_data_inst.sprite_data[125] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[126]$_DFF_PN1_  (.CLK(\clknet_5_7__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net76),
    .D(_0057_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[126] ),
    .Q(_1087_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[127]$_DFF_PN1_  (.CLK(\clknet_5_15__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net76),
    .D(_0977_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[127] ),
    .Q(_1088_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[128]$_DFF_PN0_  (.CLK(\clknet_5_15__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net76),
    .D(\top_inst.sprite_data_inst.sprite_data[129] ),
    .Q_N(_0977_),
    .Q(\top_inst.sprite_data_inst.sprite_data[128] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[129]$_DFF_PN1_  (.CLK(\clknet_5_14__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net63),
    .D(_1034_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[129] ),
    .Q(_1089_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[12]$_DFF_PN0_  (.CLK(\clknet_5_27__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net80),
    .D(\top_inst.sprite_data_inst.sprite_data[13] ),
    .Q_N(_1033_),
    .Q(\top_inst.sprite_data_inst.sprite_data[12] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[130]$_DFF_PN0_  (.CLK(\clknet_5_14__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net63),
    .D(\top_inst.sprite_data_inst.sprite_data[131] ),
    .Q_N(_1034_),
    .Q(\top_inst.sprite_data_inst.sprite_data[130] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[131]$_DFF_PN0_  (.CLK(\clknet_5_14__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net63),
    .D(\top_inst.sprite_data_inst.sprite_data[132] ),
    .Q_N(_1035_),
    .Q(\top_inst.sprite_data_inst.sprite_data[131] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[132]$_DFF_PN0_  (.CLK(\clknet_5_12__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net61),
    .D(\top_inst.sprite_data_inst.sprite_data[133] ),
    .Q_N(_1036_),
    .Q(\top_inst.sprite_data_inst.sprite_data[132] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[133]$_DFF_PN0_  (.CLK(\clknet_5_11__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net61),
    .D(\top_inst.sprite_data_inst.sprite_data[134] ),
    .Q_N(_1037_),
    .Q(\top_inst.sprite_data_inst.sprite_data[133] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[134]$_DFF_PN0_  (.CLK(\clknet_5_13__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net61),
    .D(\top_inst.sprite_data_inst.sprite_data[135] ),
    .Q_N(_0976_),
    .Q(\top_inst.sprite_data_inst.sprite_data[134] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[135]$_DFF_PN1_  (.CLK(\clknet_5_15__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net76),
    .D(_0058_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[135] ),
    .Q(_1090_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[136]$_DFF_PN1_  (.CLK(\clknet_5_24__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net76),
    .D(_0059_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[136] ),
    .Q(_1091_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[137]$_DFF_PN1_  (.CLK(\clknet_5_25__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net84),
    .D(_0060_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[137] ),
    .Q(_1092_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[138]$_DFF_PN1_  (.CLK(\clknet_5_26__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net80),
    .D(_0061_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[138] ),
    .Q(_1093_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[139]$_DFF_PN1_  (.CLK(\clknet_5_26__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net88),
    .D(_1039_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[139] ),
    .Q(_1094_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[13]$_DFF_PN0_  (.CLK(\clknet_5_24__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net80),
    .D(\top_inst.sprite_data_inst.sprite_data[14] ),
    .Q_N(_1038_),
    .Q(\top_inst.sprite_data_inst.sprite_data[13] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[140]$_DFF_PN0_  (.CLK(\clknet_5_26__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net88),
    .D(\top_inst.sprite_data_inst.sprite_data[141] ),
    .Q_N(_1039_),
    .Q(\top_inst.sprite_data_inst.sprite_data[140] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[141]$_DFF_PN0_  (.CLK(\clknet_5_28__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net88),
    .D(\top_inst.sprite_data_inst.sprite_data[142] ),
    .Q_N(_1040_),
    .Q(\top_inst.sprite_data_inst.sprite_data[141] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[142]$_DFF_PN0_  (.CLK(\clknet_5_30__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net88),
    .D(\top_inst.sprite_data_inst.sprite_data[143] ),
    .Q_N(_1041_),
    .Q(\top_inst.sprite_data_inst.sprite_data[142] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[143]$_DFF_PN0_  (.CLK(\clknet_5_26__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net88),
    .D(\top_inst.sprite_data_inst.new_sprite_data ),
    .Q_N(_0975_),
    .Q(\top_inst.sprite_data_inst.sprite_data[143] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[14]$_DFF_PN1_  (.CLK(\clknet_5_24__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net80),
    .D(_1042_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[14] ),
    .Q(_1095_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[15]$_DFF_PN0_  (.CLK(\clknet_5_24__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net81),
    .D(\top_inst.sprite_data_inst.sprite_data[16] ),
    .Q_N(_1042_),
    .Q(\top_inst.sprite_data_inst.sprite_data[15] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[16]$_DFF_PN0_  (.CLK(\clknet_5_24__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net81),
    .D(\top_inst.sprite_data_inst.sprite_data[17] ),
    .Q_N(_1043_),
    .Q(\top_inst.sprite_data_inst.sprite_data[16] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[17]$_DFF_PN0_  (.CLK(\clknet_5_15__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net81),
    .D(\top_inst.sprite_data_inst.sprite_data[18] ),
    .Q_N(_1044_),
    .Q(\top_inst.sprite_data_inst.sprite_data[17] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[18]$_DFF_PN0_  (.CLK(\clknet_5_14__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net66),
    .D(\top_inst.sprite_data_inst.sprite_data[19] ),
    .Q_N(_1045_),
    .Q(\top_inst.sprite_data_inst.sprite_data[18] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[19]$_DFF_PN0_  (.CLK(\clknet_5_14__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net66),
    .D(\top_inst.sprite_data_inst.sprite_data[20] ),
    .Q_N(_1046_),
    .Q(\top_inst.sprite_data_inst.sprite_data[19] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[1]$_DFF_PN0_  (.CLK(\clknet_5_30__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net89),
    .D(\top_inst.sprite_data_inst.sprite_data[2] ),
    .Q_N(_1047_),
    .Q(\top_inst.sprite_data_inst.sprite_data[1] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[20]$_DFF_PN0_  (.CLK(\clknet_5_13__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net66),
    .D(\top_inst.sprite_data_inst.sprite_data[21] ),
    .Q_N(_0974_),
    .Q(\top_inst.sprite_data_inst.sprite_data[20] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[21]$_DFF_PN1_  (.CLK(\clknet_5_13__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net65),
    .D(_1048_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[21] ),
    .Q(_1096_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[22]$_DFF_PN0_  (.CLK(\clknet_5_10__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net65),
    .D(\top_inst.sprite_data_inst.sprite_data[23] ),
    .Q_N(_1048_),
    .Q(\top_inst.sprite_data_inst.sprite_data[22] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[23]$_DFF_PN0_  (.CLK(\clknet_5_10__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net61),
    .D(\top_inst.sprite_data_inst.sprite_data[24] ),
    .Q_N(_1049_),
    .Q(\top_inst.sprite_data_inst.sprite_data[23] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[24]$_DFF_PN0_  (.CLK(\clknet_5_11__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net56),
    .D(\top_inst.sprite_data_inst.sprite_data[25] ),
    .Q_N(_0973_),
    .Q(\top_inst.sprite_data_inst.sprite_data[24] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[25]$_DFF_PN1_  (.CLK(\clknet_5_9__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net57),
    .D(_0062_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[25] ),
    .Q(_1097_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[26]$_DFF_PN1_  (.CLK(\clknet_5_9__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net57),
    .D(_0063_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[26] ),
    .Q(_1098_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[27]$_DFF_PN1_  (.CLK(\clknet_5_10__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net57),
    .D(_0064_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[27] ),
    .Q(_1099_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[28]$_DFF_PN1_  (.CLK(\clknet_5_13__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net61),
    .D(_0065_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[28] ),
    .Q(_1100_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[29]$_DFF_PN1_  (.CLK(\clknet_5_12__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net61),
    .D(_0066_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[29] ),
    .Q(_1101_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[2]$_DFF_PN0_  (.CLK(\clknet_5_31__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net89),
    .D(\top_inst.sprite_data_inst.sprite_data[3] ),
    .Q_N(_0972_),
    .Q(\top_inst.sprite_data_inst.sprite_data[2] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[30]$_DFF_PN1_  (.CLK(\clknet_5_12__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net60),
    .D(_1050_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[30] ),
    .Q(_1102_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[31]$_DFF_PN0_  (.CLK(\clknet_5_12__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net60),
    .D(\top_inst.sprite_data_inst.sprite_data[32] ),
    .Q_N(_1050_),
    .Q(\top_inst.sprite_data_inst.sprite_data[31] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[32]$_DFF_PN0_  (.CLK(\clknet_5_0__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net60),
    .D(\top_inst.sprite_data_inst.sprite_data[33] ),
    .Q_N(_1051_),
    .Q(\top_inst.sprite_data_inst.sprite_data[32] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[33]$_DFF_PN0_  (.CLK(\clknet_5_3__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net56),
    .D(\top_inst.sprite_data_inst.sprite_data[34] ),
    .Q_N(_0971_),
    .Q(\top_inst.sprite_data_inst.sprite_data[33] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[34]$_DFF_PN1_  (.CLK(\clknet_5_2__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net56),
    .D(_0970_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[34] ),
    .Q(_1103_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[35]$_DFF_PN0_  (.CLK(\clknet_5_2__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net56),
    .D(\top_inst.sprite_data_inst.sprite_data[36] ),
    .Q_N(_0970_),
    .Q(\top_inst.sprite_data_inst.sprite_data[35] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[36]$_DFF_PN1_  (.CLK(\clknet_5_3__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net54),
    .D(_0067_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[36] ),
    .Q(_1104_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[37]$_DFF_PN1_  (.CLK(\clknet_5_3__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net54),
    .D(_0068_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[37] ),
    .Q(_1105_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[38]$_DFF_PN1_  (.CLK(\clknet_5_2__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net54),
    .D(_0069_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[38] ),
    .Q(_1106_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[39]$_DFF_PN1_  (.CLK(\clknet_5_2__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net54),
    .D(_0070_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[39] ),
    .Q(_1107_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[3]$_DFF_PN1_  (.CLK(\clknet_5_31__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net89),
    .D(_0071_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[3] ),
    .Q(_1108_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[40]$_DFF_PN1_  (.CLK(\clknet_5_0__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net54),
    .D(_0072_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[40] ),
    .Q(_1109_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[41]$_DFF_PN1_  (.CLK(\clknet_5_0__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net56),
    .D(_0073_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[41] ),
    .Q(_1110_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[42]$_DFF_PN1_  (.CLK(\clknet_5_4__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net62),
    .D(_1052_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[42] ),
    .Q(_1111_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[43]$_DFF_PN0_  (.CLK(\clknet_5_4__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net62),
    .D(\top_inst.sprite_data_inst.sprite_data[44] ),
    .Q_N(_1052_),
    .Q(\top_inst.sprite_data_inst.sprite_data[43] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[44]$_DFF_PN0_  (.CLK(\clknet_5_4__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net60),
    .D(\top_inst.sprite_data_inst.sprite_data[45] ),
    .Q_N(_1053_),
    .Q(\top_inst.sprite_data_inst.sprite_data[44] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[45]$_DFF_PN0_  (.CLK(\clknet_5_1__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net60),
    .D(\top_inst.sprite_data_inst.sprite_data[46] ),
    .Q_N(_1054_),
    .Q(\top_inst.sprite_data_inst.sprite_data[45] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[46]$_DFF_PN0_  (.CLK(\clknet_5_1__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net60),
    .D(\top_inst.sprite_data_inst.sprite_data[47] ),
    .Q_N(_0969_),
    .Q(\top_inst.sprite_data_inst.sprite_data[46] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[47]$_DFF_PN1_  (.CLK(\clknet_5_1__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net56),
    .D(_1055_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[47] ),
    .Q(_1112_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[48]$_DFF_PN0_  (.CLK(\clknet_5_0__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net56),
    .D(\top_inst.sprite_data_inst.sprite_data[49] ),
    .Q_N(_1055_),
    .Q(\top_inst.sprite_data_inst.sprite_data[48] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[49]$_DFF_PN0_  (.CLK(\clknet_5_0__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net56),
    .D(\top_inst.sprite_data_inst.sprite_data[50] ),
    .Q_N(_0968_),
    .Q(\top_inst.sprite_data_inst.sprite_data[49] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[4]$_DFF_PN1_  (.CLK(\clknet_5_31__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net90),
    .D(_0074_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[4] ),
    .Q(_1113_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[50]$_DFF_PN0_  (.CLK(\clknet_5_3__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net54),
    .D(\top_inst.sprite_data_inst.sprite_data[51] ),
    .Q_N(_0967_),
    .Q(\top_inst.sprite_data_inst.sprite_data[50] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[51]$_DFF_PN1_  (.CLK(\clknet_5_2__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net54),
    .D(_0075_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[51] ),
    .Q(_1114_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[52]$_DFF_PN1_  (.CLK(\clknet_5_11__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net60),
    .D(_1056_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[52] ),
    .Q(_1115_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[53]$_DFF_PN0_  (.CLK(\clknet_5_12__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net64),
    .D(\top_inst.sprite_data_inst.sprite_data[54] ),
    .Q_N(_1056_),
    .Q(\top_inst.sprite_data_inst.sprite_data[53] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[54]$_DFF_PN0_  (.CLK(\clknet_5_11__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net64),
    .D(\top_inst.sprite_data_inst.sprite_data[55] ),
    .Q_N(_1057_),
    .Q(\top_inst.sprite_data_inst.sprite_data[54] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[55]$_DFF_PN0_  (.CLK(\clknet_5_10__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net57),
    .D(\top_inst.sprite_data_inst.sprite_data[56] ),
    .Q_N(_1058_),
    .Q(\top_inst.sprite_data_inst.sprite_data[55] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[56]$_DFF_PN0_  (.CLK(\clknet_5_9__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net57),
    .D(\top_inst.sprite_data_inst.sprite_data[57] ),
    .Q_N(_1059_),
    .Q(\top_inst.sprite_data_inst.sprite_data[56] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[57]$_DFF_PN0_  (.CLK(\clknet_5_8__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net54),
    .D(\top_inst.sprite_data_inst.sprite_data[58] ),
    .Q_N(_1060_),
    .Q(\top_inst.sprite_data_inst.sprite_data[57] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[58]$_DFF_PN0_  (.CLK(\clknet_5_8__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net55),
    .D(\top_inst.sprite_data_inst.sprite_data[59] ),
    .Q_N(_0966_),
    .Q(\top_inst.sprite_data_inst.sprite_data[58] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[59]$_DFF_PN1_  (.CLK(\clknet_5_8__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net55),
    .D(_0076_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[59] ),
    .Q(_1116_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[5]$_DFF_PN1_  (.CLK(\clknet_5_30__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net90),
    .D(_0077_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[5] ),
    .Q(_1117_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[60]$_DFF_PN1_  (.CLK(\clknet_5_9__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net55),
    .D(_1061_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[60] ),
    .Q(_1118_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[61]$_DFF_PN0_  (.CLK(\clknet_5_8__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net55),
    .D(\top_inst.sprite_data_inst.sprite_data[62] ),
    .Q_N(_1061_),
    .Q(\top_inst.sprite_data_inst.sprite_data[61] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[62]$_DFF_PN0_  (.CLK(\clknet_5_8__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net55),
    .D(\top_inst.sprite_data_inst.sprite_data[63] ),
    .Q_N(_0965_),
    .Q(\top_inst.sprite_data_inst.sprite_data[62] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[63]$_DFF_PN1_  (.CLK(\clknet_5_10__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net57),
    .D(_0078_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[63] ),
    .Q(_1119_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[64]$_DFF_PN1_  (.CLK(\clknet_5_6__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net63),
    .D(_0079_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[64] ),
    .Q(_1120_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[65]$_DFF_PN1_  (.CLK(\clknet_5_6__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net63),
    .D(_0080_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[65] ),
    .Q(_1121_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[66]$_DFF_PN1_  (.CLK(\clknet_5_6__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net62),
    .D(_0081_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[66] ),
    .Q(_1122_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[67]$_DFF_PN1_  (.CLK(\clknet_5_5__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net62),
    .D(_0082_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[67] ),
    .Q(_1123_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[68]$_DFF_PN1_  (.CLK(\clknet_5_6__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net62),
    .D(_0083_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[68] ),
    .Q(_1124_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[69]$_DFF_PN1_  (.CLK(\clknet_5_4__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net61),
    .D(_0964_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[69] ),
    .Q(_1125_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[6]$_DFF_PN1_  (.CLK(\clknet_5_30__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net89),
    .D(_0084_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[6] ),
    .Q(_1126_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[70]$_DFF_PN0_  (.CLK(\clknet_5_1__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net60),
    .D(\top_inst.sprite_data_inst.sprite_data[71] ),
    .Q_N(_0964_),
    .Q(\top_inst.sprite_data_inst.sprite_data[70] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[71]$_DFF_PN1_  (.CLK(\clknet_5_4__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net62),
    .D(_0085_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[71] ),
    .Q(_1127_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[72]$_DFF_PN1_  (.CLK(\clknet_5_5__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net75),
    .D(_1062_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[72] ),
    .Q(_1128_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[73]$_DFF_PN0_  (.CLK(\clknet_5_17__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net77),
    .D(\top_inst.sprite_data_inst.sprite_data[74] ),
    .Q_N(_1062_),
    .Q(\top_inst.sprite_data_inst.sprite_data[73] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[74]$_DFF_PN0_  (.CLK(\clknet_5_16__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net75),
    .D(\top_inst.sprite_data_inst.sprite_data[75] ),
    .Q_N(_0963_),
    .Q(\top_inst.sprite_data_inst.sprite_data[74] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[75]$_DFF_PN1_  (.CLK(\clknet_5_5__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net75),
    .D(_0086_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[75] ),
    .Q(_1129_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[76]$_DFF_PN1_  (.CLK(\clknet_5_7__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net75),
    .D(_0087_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[76] ),
    .Q(_1130_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[77]$_DFF_PN1_  (.CLK(\clknet_5_5__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net62),
    .D(_0088_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[77] ),
    .Q(_1131_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[78]$_DFF_PN1_  (.CLK(\clknet_5_6__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net62),
    .D(_0089_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[78] ),
    .Q(_1132_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[79]$_DFF_PN1_  (.CLK(\clknet_5_18__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net78),
    .D(_0090_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[79] ),
    .Q(_1133_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[7]$_DFF_PN1_  (.CLK(\clknet_5_30__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net89),
    .D(_0091_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[7] ),
    .Q(_1134_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[80]$_DFF_PN1_  (.CLK(\clknet_5_18__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net78),
    .D(_0092_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[80] ),
    .Q(_1135_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[81]$_DFF_PN1_  (.CLK(\clknet_5_25__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net78),
    .D(_0962_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[81] ),
    .Q(_1136_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[82]$_DFF_PN0_  (.CLK(\clknet_5_25__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net78),
    .D(\top_inst.sprite_data_inst.sprite_data[83] ),
    .Q_N(_0962_),
    .Q(\top_inst.sprite_data_inst.sprite_data[82] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[83]$_DFF_PN1_  (.CLK(\clknet_5_25__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net78),
    .D(_0093_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[83] ),
    .Q(_1137_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[84]$_DFF_PN1_  (.CLK(\clknet_5_27__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net84),
    .D(_1063_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[84] ),
    .Q(_1138_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[85]$_DFF_PN0_  (.CLK(\clknet_5_29__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net85),
    .D(\top_inst.sprite_data_inst.sprite_data[86] ),
    .Q_N(_1063_),
    .Q(\top_inst.sprite_data_inst.sprite_data[85] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[86]$_DFF_PN0_  (.CLK(\clknet_5_28__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net84),
    .D(\top_inst.sprite_data_inst.sprite_data[87] ),
    .Q_N(_0961_),
    .Q(\top_inst.sprite_data_inst.sprite_data[86] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[87]$_DFF_PN1_  (.CLK(\clknet_5_28__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net84),
    .D(_0094_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[87] ),
    .Q(_1139_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[88]$_DFF_PN1_  (.CLK(\clknet_5_29__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net85),
    .D(_0960_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[88] ),
    .Q(_1140_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[89]$_DFF_PN0_  (.CLK(\clknet_5_29__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net86),
    .D(\top_inst.sprite_data_inst.sprite_data[90] ),
    .Q_N(_0960_),
    .Q(\top_inst.sprite_data_inst.sprite_data[89] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[8]$_DFF_PN1_  (.CLK(\clknet_5_29__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net89),
    .D(_0957_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[8] ),
    .Q(_1141_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[90]$_DFF_PN1_  (.CLK(\clknet_5_28__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net86),
    .D(_0095_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[90] ),
    .Q(_1142_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[91]$_DFF_PN1_  (.CLK(\clknet_5_22__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net84),
    .D(_1064_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[91] ),
    .Q(_1143_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[92]$_DFF_PN0_  (.CLK(\clknet_5_27__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net84),
    .D(\top_inst.sprite_data_inst.sprite_data[93] ),
    .Q_N(_1064_),
    .Q(\top_inst.sprite_data_inst.sprite_data[92] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[93]$_DFF_PN0_  (.CLK(\clknet_5_22__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net87),
    .D(\top_inst.sprite_data_inst.sprite_data[94] ),
    .Q_N(_1065_),
    .Q(\top_inst.sprite_data_inst.sprite_data[93] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[94]$_DFF_PN0_  (.CLK(\clknet_5_18__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net78),
    .D(\top_inst.sprite_data_inst.sprite_data[95] ),
    .Q_N(_0959_),
    .Q(\top_inst.sprite_data_inst.sprite_data[94] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[95]$_DFF_PN1_  (.CLK(\clknet_5_19__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net79),
    .D(_0096_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[95] ),
    .Q(_1144_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[96]$_DFF_PN1_  (.CLK(\clknet_5_23__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net86),
    .D(_1066_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[96] ),
    .Q(_1145_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[97]$_DFF_PN0_  (.CLK(\clknet_5_20__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net86),
    .D(\top_inst.sprite_data_inst.sprite_data[98] ),
    .Q_N(_1066_),
    .Q(\top_inst.sprite_data_inst.sprite_data[97] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[98]$_DFF_PN0_  (.CLK(\clknet_5_22__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net84),
    .D(\top_inst.sprite_data_inst.sprite_data[99] ),
    .Q_N(_0958_),
    .Q(\top_inst.sprite_data_inst.sprite_data[98] ));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[99]$_DFF_PN1_  (.CLK(\clknet_5_22__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net83),
    .D(_0097_),
    .Q_N(\top_inst.sprite_data_inst.sprite_data[99] ),
    .Q(_1146_));
 sg13g2_dfrbp_1 \top_inst.sprite_data_inst.sprite_data[9]$_DFF_PN0_  (.CLK(\clknet_5_28__leaf_top_inst.sprite_data_inst.gclk ),
    .RESET_B(net89),
    .D(\top_inst.sprite_data_inst.sprite_data[10] ),
    .Q_N(_0957_),
    .Q(\top_inst.sprite_data_inst.sprite_data[9] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.divider$_DFFE_PN0P_  (.CLK(clknet_level_3_1_1351_clk),
    .RESET_B(net72),
    .D(_0139_),
    .Q_N(_0029_),
    .Q(\top_inst.sprite_movement_inst.divider ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_x[0]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_13_clk),
    .RESET_B(net67),
    .D(_0140_),
    .Q_N(_0045_),
    .Q(\top_inst.sprite_movement_inst.sprite_x[0] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_x[1]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_13_clk),
    .RESET_B(net59),
    .D(_0141_),
    .Q_N(_0956_),
    .Q(\top_inst.sprite_movement_inst.sprite_x[1] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_x[2]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_13_clk),
    .RESET_B(net59),
    .D(_0142_),
    .Q_N(_0955_),
    .Q(\top_inst.sprite_movement_inst.sprite_x[2] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_x[3]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_13_clk),
    .RESET_B(net59),
    .D(_0143_),
    .Q_N(_0954_),
    .Q(\top_inst.sprite_movement_inst.sprite_x[3] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_x[4]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_311_clk),
    .RESET_B(net59),
    .D(_0144_),
    .Q_N(_0953_),
    .Q(\top_inst.sprite_movement_inst.sprite_x[4] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_x[5]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_13_clk),
    .RESET_B(net67),
    .D(_0145_),
    .Q_N(_0952_),
    .Q(\top_inst.sprite_movement_inst.sprite_x[5] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_x[6]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_13_clk),
    .RESET_B(net67),
    .D(_0146_),
    .Q_N(_0951_),
    .Q(\top_inst.sprite_movement_inst.sprite_x[6] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_x[7]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_27_clk),
    .RESET_B(net67),
    .D(_0147_),
    .Q_N(_0950_),
    .Q(\top_inst.sprite_movement_inst.sprite_x[7] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_x_dir$_DFFE_PN0P_  (.CLK(clknet_level_3_1_13_clk),
    .RESET_B(net59),
    .D(_0148_),
    .Q_N(_0949_),
    .Q(\top_inst.sprite_movement_inst.sprite_x_dir ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_y[0]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_27_clk),
    .RESET_B(net67),
    .D(_0149_),
    .Q_N(_0046_),
    .Q(\top_inst.sprite_movement_inst.sprite_y[0] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_y[1]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_27_clk),
    .RESET_B(net67),
    .D(_0150_),
    .Q_N(_0948_),
    .Q(\top_inst.sprite_movement_inst.sprite_y[1] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_y[2]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_27_clk),
    .RESET_B(net71),
    .D(_0151_),
    .Q_N(_0947_),
    .Q(\top_inst.sprite_movement_inst.sprite_y[2] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_y[3]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_27_clk),
    .RESET_B(net71),
    .D(_0152_),
    .Q_N(_0946_),
    .Q(\top_inst.sprite_movement_inst.sprite_y[3] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_y[4]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_519_clk),
    .RESET_B(net71),
    .D(_0153_),
    .Q_N(_0945_),
    .Q(\top_inst.sprite_movement_inst.sprite_y[4] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_y[5]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_519_clk),
    .RESET_B(net68),
    .D(_0154_),
    .Q_N(_0944_),
    .Q(\top_inst.sprite_movement_inst.sprite_y[5] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_y[6]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_519_clk),
    .RESET_B(net67),
    .D(_0155_),
    .Q_N(_0943_),
    .Q(\top_inst.sprite_movement_inst.sprite_y[6] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_y[7]$_DFFE_PN0P_  (.CLK(clknet_level_3_1_519_clk),
    .RESET_B(net68),
    .D(_0156_),
    .Q_N(_0942_),
    .Q(\top_inst.sprite_movement_inst.sprite_y[7] ));
 sg13g2_dfrbp_1 \top_inst.sprite_movement_inst.sprite_y_dir$_DFFE_PN0P_  (.CLK(clknet_level_3_1_27_clk),
    .RESET_B(net67),
    .D(_0157_),
    .Q_N(_0941_),
    .Q(\top_inst.sprite_movement_inst.sprite_y_dir ));
 sg13g2_dfrbp_1 \top_inst.sprite_x[0]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_415_clk),
    .RESET_B(net65),
    .D(_0158_),
    .Q_N(_0940_),
    .Q(\top_inst.sprite_x[0] ));
 sg13g2_dfrbp_1 \top_inst.sprite_x[1]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_311_clk),
    .RESET_B(net65),
    .D(_0159_),
    .Q_N(_0939_),
    .Q(\top_inst.sprite_x[1] ));
 sg13g2_dfrbp_1 \top_inst.sprite_x[2]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_311_clk),
    .RESET_B(net59),
    .D(_0160_),
    .Q_N(_0938_),
    .Q(\top_inst.sprite_x[2] ));
 sg13g2_dfrbp_1 \top_inst.sprite_x[3]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_311_clk),
    .RESET_B(net65),
    .D(_0161_),
    .Q_N(_0937_),
    .Q(\top_inst.sprite_x[3] ));
 sg13g2_dfrbp_1 \top_inst.sprite_x[4]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_415_clk),
    .RESET_B(net66),
    .D(_0162_),
    .Q_N(_0936_),
    .Q(\top_inst.sprite_x[4] ));
 sg13g2_dfrbp_1 \top_inst.sprite_x[5]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_311_clk),
    .RESET_B(net65),
    .D(_0163_),
    .Q_N(_0935_),
    .Q(\top_inst.sprite_x[5] ));
 sg13g2_dfrbp_1 \top_inst.sprite_x[6]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_311_clk),
    .RESET_B(net65),
    .D(_0164_),
    .Q_N(_0934_),
    .Q(\top_inst.sprite_x[6] ));
 sg13g2_dfrbp_1 \top_inst.sprite_x[7]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_311_clk),
    .RESET_B(net65),
    .D(_0165_),
    .Q_N(_0933_),
    .Q(\top_inst.sprite_x[7] ));
 sg13g2_dfrbp_1 \top_inst.sprite_y[0]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_727_clk),
    .RESET_B(net72),
    .D(_0166_),
    .Q_N(_0932_),
    .Q(\top_inst.sprite_y[0] ));
 sg13g2_dfrbp_1 \top_inst.sprite_y[1]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_1351_clk),
    .RESET_B(net72),
    .D(_0167_),
    .Q_N(_0931_),
    .Q(\top_inst.sprite_y[1] ));
 sg13g2_dfrbp_1 \top_inst.sprite_y[2]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_415_clk),
    .RESET_B(net72),
    .D(_0168_),
    .Q_N(_0930_),
    .Q(\top_inst.sprite_y[2] ));
 sg13g2_dfrbp_1 \top_inst.sprite_y[3]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_415_clk),
    .RESET_B(net72),
    .D(_0169_),
    .Q_N(_0929_),
    .Q(\top_inst.sprite_y[3] ));
 sg13g2_dfrbp_1 \top_inst.sprite_y[4]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_27_clk),
    .RESET_B(net72),
    .D(_0170_),
    .Q_N(_0928_),
    .Q(\top_inst.sprite_y[4] ));
 sg13g2_dfrbp_1 \top_inst.sprite_y[5]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_415_clk),
    .RESET_B(net72),
    .D(_0171_),
    .Q_N(_0927_),
    .Q(\top_inst.sprite_y[5] ));
 sg13g2_dfrbp_1 \top_inst.sprite_y[6]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_415_clk),
    .RESET_B(net72),
    .D(_0172_),
    .Q_N(_0926_),
    .Q(\top_inst.sprite_y[6] ));
 sg13g2_dfrbp_1 \top_inst.sprite_y[7]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_415_clk),
    .RESET_B(net66),
    .D(_0173_),
    .Q_N(_1067_),
    .Q(\top_inst.sprite_y[7] ));
 sg13g2_dfrbp_1 \top_inst.synchronizer_spi_cs.pipe[0]$_DFF_PN0_  (.CLK(clknet_level_3_1_1663_clk),
    .RESET_B(net93),
    .D(net3),
    .Q_N(_1068_),
    .Q(\top_inst.synchronizer_spi_cs.pipe[0] ));
 sg13g2_dfrbp_1 \top_inst.synchronizer_spi_cs.pipe[1]$_DFF_PN0_  (.CLK(clknet_level_3_1_1663_clk),
    .RESET_B(net93),
    .D(\top_inst.synchronizer_spi_cs.pipe[0] ),
    .Q_N(_1069_),
    .Q(\top_inst.spi_cs_sync ));
 sg13g2_dfrbp_1 \top_inst.synchronizer_spi_mosi.pipe[0]$_DFF_PN0_  (.CLK(clknet_level_3_1_1455_clk),
    .RESET_B(net94),
    .D(net4),
    .Q_N(_1070_),
    .Q(\top_inst.synchronizer_spi_mosi.pipe[0] ));
 sg13g2_dfrbp_1 \top_inst.synchronizer_spi_mosi.pipe[1]$_DFF_PN0_  (.CLK(clknet_level_3_1_1351_clk),
    .RESET_B(net94),
    .D(\top_inst.synchronizer_spi_mosi.pipe[0] ),
    .Q_N(_1071_),
    .Q(\top_inst.spi_mosi_sync ));
 sg13g2_dfrbp_1 \top_inst.synchronizer_spi_sclk.pipe[0]$_DFF_PN0_  (.CLK(clknet_level_3_1_1351_clk),
    .RESET_B(net94),
    .D(net5),
    .Q_N(_1072_),
    .Q(\top_inst.synchronizer_spi_sclk.pipe[0] ));
 sg13g2_dfrbp_1 \top_inst.synchronizer_spi_sclk.pipe[1]$_DFF_PN0_  (.CLK(clknet_level_3_1_1455_clk),
    .RESET_B(net93),
    .D(\top_inst.synchronizer_spi_sclk.pipe[0] ),
    .Q_N(_0925_),
    .Q(\top_inst.spi_receiver_inst.spi_sclk ));
 sg13g2_dfrbp_1 \top_inst.time_dir$_DFFE_PN0P_  (.CLK(clknet_level_3_1_1247_clk),
    .RESET_B(net92),
    .D(_0174_),
    .Q_N(_1073_),
    .Q(\top_inst.time_dir ));
 sg13g2_dfrbp_1 \top_inst.timing_hor.counter[0]$_DFF_PN0_  (.CLK(clknet_level_3_1_1143_clk),
    .RESET_B(net88),
    .D(_0030_),
    .Q_N(_0924_),
    .Q(\top_inst.background_inst.counter_h[0] ));
 sg13g2_dfrbp_1 \top_inst.timing_hor.counter[10]$_DFF_PN1_  (.CLK(clknet_level_3_1_935_clk),
    .RESET_B(net80),
    .D(_0098_),
    .Q_N(\top_inst.background_inst.counter_h[10] ),
    .Q(_1147_));
 sg13g2_dfrbp_1 \top_inst.timing_hor.counter[11]$_DFF_PN1_  (.CLK(clknet_level_3_1_935_clk),
    .RESET_B(net80),
    .D(_0099_),
    .Q_N(\top_inst.background_inst.counter_h[11] ),
    .Q(_1148_));
 sg13g2_dfrbp_1 \top_inst.timing_hor.counter[1]$_DFF_PN0_  (.CLK(clknet_level_3_1_1143_clk),
    .RESET_B(net90),
    .D(_0031_),
    .Q_N(_1074_),
    .Q(\top_inst.background_inst.counter_h[1] ));
 sg13g2_dfrbp_1 \top_inst.timing_hor.counter[2]$_DFF_PN0_  (.CLK(clknet_level_3_1_1247_clk),
    .RESET_B(net90),
    .D(_0032_),
    .Q_N(_1075_),
    .Q(\top_inst.background_inst.counter_h[2] ));
 sg13g2_dfrbp_1 \top_inst.timing_hor.counter[3]$_DFF_PN0_  (.CLK(clknet_level_3_1_1143_clk),
    .RESET_B(net90),
    .D(_0033_),
    .Q_N(_1076_),
    .Q(\top_inst.background_inst.counter_h[3] ));
 sg13g2_dfrbp_1 \top_inst.timing_hor.counter[4]$_DFF_PN0_  (.CLK(clknet_level_3_1_1143_clk),
    .RESET_B(net80),
    .D(_0034_),
    .Q_N(_1077_),
    .Q(\top_inst.background_inst.counter_h[4] ));
 sg13g2_dfrbp_1 \top_inst.timing_hor.counter[5]$_DFF_PN0_  (.CLK(clknet_level_3_1_935_clk),
    .RESET_B(net82),
    .D(_0035_),
    .Q_N(_0038_),
    .Q(\top_inst.background_inst.counter_h[5] ));
 sg13g2_dfrbp_1 \top_inst.timing_hor.counter[6]$_DFF_PN0_  (.CLK(clknet_level_3_1_1039_clk),
    .RESET_B(net81),
    .D(_0036_),
    .Q_N(_0040_),
    .Q(\top_inst.background_inst.counter_h[6] ));
 sg13g2_dfrbp_1 \top_inst.timing_hor.counter[7]$_DFF_PN0_  (.CLK(clknet_level_3_1_935_clk),
    .RESET_B(net81),
    .D(_0037_),
    .Q_N(_0923_),
    .Q(\top_inst.background_inst.counter_h[7] ));
 sg13g2_dfrbp_1 \top_inst.timing_hor.counter[8]$_DFF_PN1_  (.CLK(clknet_level_3_1_935_clk),
    .RESET_B(net81),
    .D(_0100_),
    .Q_N(\top_inst.background_inst.counter_h[8] ),
    .Q(_1149_));
 sg13g2_dfrbp_1 \top_inst.timing_hor.counter[9]$_DFF_PN1_  (.CLK(clknet_level_3_1_935_clk),
    .RESET_B(net80),
    .D(_0101_),
    .Q_N(\top_inst.background_inst.counter_h[9] ),
    .Q(_1150_));
 sg13g2_dfrbp_1 \top_inst.timing_ver.counter[0]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_1351_clk),
    .RESET_B(net91),
    .D(_0175_),
    .Q_N(_0042_),
    .Q(\top_inst.background_inst.counter_v[0] ));
 sg13g2_dfrbp_1 \top_inst.timing_ver.counter[10]$_DFFE_PN1N_  (.CLK(clknet_level_3_1_1039_clk),
    .RESET_B(net81),
    .D(_0176_),
    .Q_N(\top_inst.background_inst.counter_v[10] ),
    .Q(_0048_));
 sg13g2_dfrbp_1 \top_inst.timing_ver.counter[1]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_1247_clk),
    .RESET_B(net92),
    .D(_0177_),
    .Q_N(_0922_),
    .Q(\top_inst.background_inst.counter_v[1] ));
 sg13g2_dfrbp_1 \top_inst.timing_ver.counter[2]$_DFFE_PN1N_  (.CLK(clknet_level_3_1_1143_clk),
    .RESET_B(net82),
    .D(_0178_),
    .Q_N(\top_inst.background_inst.counter_v[2] ),
    .Q(_0049_));
 sg13g2_dfrbp_1 \top_inst.timing_ver.counter[3]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_1143_clk),
    .RESET_B(net91),
    .D(_0179_),
    .Q_N(_0039_),
    .Q(\top_inst.background_inst.counter_v[3] ));
 sg13g2_dfrbp_1 \top_inst.timing_ver.counter[4]$_DFFE_PN0N_  (.CLK(clknet_level_3_1_1039_clk),
    .RESET_B(net91),
    .D(_0180_),
    .Q_N(_0921_),
    .Q(\top_inst.background_inst.counter_v[4] ));
 sg13g2_dfrbp_1 \top_inst.timing_ver.counter[5]$_DFFE_PN1N_  (.CLK(clknet_level_3_1_1039_clk),
    .RESET_B(net91),
    .D(_0181_),
    .Q_N(\top_inst.background_inst.counter_v[5] ),
    .Q(_0050_));
 sg13g2_dfrbp_1 \top_inst.timing_ver.counter[6]$_DFFE_PN1N_  (.CLK(clknet_level_3_1_935_clk),
    .RESET_B(net91),
    .D(_0182_),
    .Q_N(\top_inst.background_inst.counter_v[6] ),
    .Q(_0051_));
 sg13g2_dfrbp_1 \top_inst.timing_ver.counter[7]$_DFFE_PN1N_  (.CLK(clknet_level_3_1_1039_clk),
    .RESET_B(net91),
    .D(_0183_),
    .Q_N(\top_inst.background_inst.counter_v[7] ),
    .Q(_0052_));
 sg13g2_dfrbp_1 \top_inst.timing_ver.counter[8]$_DFFE_PN1N_  (.CLK(clknet_level_3_1_1039_clk),
    .RESET_B(net73),
    .D(_0184_),
    .Q_N(\top_inst.background_inst.counter_v[8] ),
    .Q(_0053_));
 sg13g2_dfrbp_1 \top_inst.timing_ver.counter[9]$_DFFE_PN1N_  (.CLK(clknet_level_3_1_1039_clk),
    .RESET_B(net91),
    .D(_0185_),
    .Q_N(\top_inst.background_inst.counter_v[9] ),
    .Q(_0054_));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(uio_in[0]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[1]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[3]),
    .X(net5));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[4]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[5]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[0]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[1]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[2]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[3]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[4]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[5]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[6]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout16 (.A(_0744_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0743_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0733_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(next_frame),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0886_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0858_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0534_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(next_vertical),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0523_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0834_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0739_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0846_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0837_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0240_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0889_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0735_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0734_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0572_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0549_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0496_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0494_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0762_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0756_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0660_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0577_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0565_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0559_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0555_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0548_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0528_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0505_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0497_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0488_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0484_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0475_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0473_),
    .X(net51));
 sg13g2_buf_1 fanout52 (.A(_0541_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0540_),
    .X(net53));
 sg13g2_buf_4 fanout54 (.X(net54),
    .A(net58));
 sg13g2_buf_2 fanout55 (.A(net58),
    .X(net55));
 sg13g2_buf_4 fanout56 (.X(net56),
    .A(net58));
 sg13g2_buf_2 fanout57 (.A(net58),
    .X(net57));
 sg13g2_buf_1 fanout58 (.A(net59),
    .X(net58));
 sg13g2_buf_4 fanout59 (.X(net59),
    .A(net74));
 sg13g2_buf_4 fanout60 (.X(net60),
    .A(net61));
 sg13g2_buf_4 fanout61 (.X(net61),
    .A(net64));
 sg13g2_buf_4 fanout62 (.X(net62),
    .A(net64));
 sg13g2_buf_2 fanout63 (.A(net64),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(net74),
    .X(net64));
 sg13g2_buf_4 fanout65 (.X(net65),
    .A(net66));
 sg13g2_buf_2 fanout66 (.A(net74),
    .X(net66));
 sg13g2_buf_4 fanout67 (.X(net67),
    .A(net71));
 sg13g2_buf_4 fanout68 (.X(net68),
    .A(net70));
 sg13g2_buf_2 fanout69 (.A(net70),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(net71),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(net74),
    .X(net71));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(net73));
 sg13g2_buf_2 fanout73 (.A(net74),
    .X(net73));
 sg13g2_buf_1 fanout74 (.A(net1),
    .X(net74));
 sg13g2_buf_4 fanout75 (.X(net75),
    .A(net79));
 sg13g2_buf_2 fanout76 (.A(net79),
    .X(net76));
 sg13g2_buf_4 fanout77 (.X(net77),
    .A(net78));
 sg13g2_buf_4 fanout78 (.X(net78),
    .A(net79));
 sg13g2_buf_1 fanout79 (.A(net82),
    .X(net79));
 sg13g2_buf_4 fanout80 (.X(net80),
    .A(net81));
 sg13g2_buf_4 fanout81 (.X(net81),
    .A(net82));
 sg13g2_buf_1 fanout82 (.A(net95),
    .X(net82));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(net84));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(net87));
 sg13g2_buf_4 fanout85 (.X(net85),
    .A(net87));
 sg13g2_buf_2 fanout86 (.A(net87),
    .X(net86));
 sg13g2_buf_1 fanout87 (.A(net95),
    .X(net87));
 sg13g2_buf_4 fanout88 (.X(net88),
    .A(net90));
 sg13g2_buf_4 fanout89 (.X(net89),
    .A(net90));
 sg13g2_buf_4 fanout90 (.X(net90),
    .A(net95));
 sg13g2_buf_4 fanout91 (.X(net91),
    .A(net94));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(net94));
 sg13g2_buf_2 fanout93 (.A(net94),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(net95),
    .X(net94));
 sg13g2_buf_1 fanout95 (.A(net1),
    .X(net95));
 sg13g2_tielo _2070__96 (.L_LO(net96));
 sg13g2_tielo _2071__97 (.L_LO(net97));
 sg13g2_tielo _2073__98 (.L_LO(net98));
 sg13g2_tielo _2076__99 (.L_LO(net99));
 sg13g2_tielo _2077__100 (.L_LO(net100));
 sg13g2_tielo _2078__101 (.L_LO(net101));
 sg13g2_tielo _2079__102 (.L_LO(net102));
 sg13g2_tielo _2080__103 (.L_LO(net103));
 sg13g2_tielo _2081__104 (.L_LO(net104));
 sg13g2_tielo _2084__105 (.L_LO(net105));
 sg13g2_tielo _2085__106 (.L_LO(net106));
 sg13g2_tiehi _2074__108 (.L_HI(net108));
 sg13g2_tiehi _2075__109 (.L_HI(net109));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[0][0]$_DLATCH_N_._TECHMAP_DLATCH_N_110  (.L_HI(net110));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[0][1]$_DLATCH_N_._TECHMAP_DLATCH_N_111  (.L_HI(net111));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[0][2]$_DLATCH_N_._TECHMAP_DLATCH_N_112  (.L_HI(net112));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[0][3]$_DLATCH_N_._TECHMAP_DLATCH_N_113  (.L_HI(net113));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[0][4]$_DLATCH_N_._TECHMAP_DLATCH_N_114  (.L_HI(net114));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[0][5]$_DLATCH_N_._TECHMAP_DLATCH_N_115  (.L_HI(net115));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[1][0]$_DLATCH_N_._TECHMAP_DLATCH_N_116  (.L_HI(net116));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[1][1]$_DLATCH_N_._TECHMAP_DLATCH_N_117  (.L_HI(net117));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[1][2]$_DLATCH_N_._TECHMAP_DLATCH_N_118  (.L_HI(net118));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[1][3]$_DLATCH_N_._TECHMAP_DLATCH_N_119  (.L_HI(net119));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[1][4]$_DLATCH_N_._TECHMAP_DLATCH_N_120  (.L_HI(net120));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[1][5]$_DLATCH_N_._TECHMAP_DLATCH_N_121  (.L_HI(net121));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[2][0]$_DLATCH_N_._TECHMAP_DLATCH_N_122  (.L_HI(net122));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[2][1]$_DLATCH_N_._TECHMAP_DLATCH_N_123  (.L_HI(net123));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[2][2]$_DLATCH_N_._TECHMAP_DLATCH_N_124  (.L_HI(net124));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[2][3]$_DLATCH_N_._TECHMAP_DLATCH_N_125  (.L_HI(net125));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[2][4]$_DLATCH_N_._TECHMAP_DLATCH_N_126  (.L_HI(net126));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[2][5]$_DLATCH_N_._TECHMAP_DLATCH_N_127  (.L_HI(net127));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[3][0]$_DLATCH_N_._TECHMAP_DLATCH_N_128  (.L_HI(net128));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[3][1]$_DLATCH_N_._TECHMAP_DLATCH_N_129  (.L_HI(net129));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[3][2]$_DLATCH_N_._TECHMAP_DLATCH_N_130  (.L_HI(net130));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[3][3]$_DLATCH_N_._TECHMAP_DLATCH_N_131  (.L_HI(net131));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[3][4]$_DLATCH_N_._TECHMAP_DLATCH_N_132  (.L_HI(net132));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[3][5]$_DLATCH_N_._TECHMAP_DLATCH_N_133  (.L_HI(net133));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[4][0]$_DLATCH_N_._TECHMAP_DLATCH_N_134  (.L_HI(net134));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[4][1]$_DLATCH_N_._TECHMAP_DLATCH_N_135  (.L_HI(net135));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[4][2]$_DLATCH_N_._TECHMAP_DLATCH_N_136  (.L_HI(net136));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[4][3]$_DLATCH_N_._TECHMAP_DLATCH_N_137  (.L_HI(net137));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[4][4]$_DLATCH_N_._TECHMAP_DLATCH_N_138  (.L_HI(net138));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[4][5]$_DLATCH_N_._TECHMAP_DLATCH_N_139  (.L_HI(net139));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[4][6]$_DLATCH_N_._TECHMAP_DLATCH_N_140  (.L_HI(net140));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[4][7]$_DLATCH_N_._TECHMAP_DLATCH_N_141  (.L_HI(net141));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[5][0]$_DLATCH_N_._TECHMAP_DLATCH_N_142  (.L_HI(net142));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[5][1]$_DLATCH_N_._TECHMAP_DLATCH_N_143  (.L_HI(net143));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[5][2]$_DLATCH_N_._TECHMAP_DLATCH_N_144  (.L_HI(net144));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[5][3]$_DLATCH_N_._TECHMAP_DLATCH_N_145  (.L_HI(net145));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[5][4]$_DLATCH_N_._TECHMAP_DLATCH_N_146  (.L_HI(net146));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[5][5]$_DLATCH_N_._TECHMAP_DLATCH_N_147  (.L_HI(net147));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[5][6]$_DLATCH_N_._TECHMAP_DLATCH_N_148  (.L_HI(net148));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[5][7]$_DLATCH_N_._TECHMAP_DLATCH_N_149  (.L_HI(net149));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[6][0]$_DLATCH_N_._TECHMAP_DLATCH_N_150  (.L_HI(net150));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[6][1]$_DLATCH_N_._TECHMAP_DLATCH_N_151  (.L_HI(net151));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[6][2]$_DLATCH_N_._TECHMAP_DLATCH_N_152  (.L_HI(net152));
 sg13g2_tiehi \top_inst.spi_receiver_inst.registers[6][3]$_DLATCH_N_._TECHMAP_DLATCH_N_153  (.L_HI(net153));
 sg13g2_tiehi \top_inst.spi_sclk_delayed$_DFF_P__154  (.L_HI(net154));
 sg13g2_tiehi \top_inst.sprite_access_inst.sprite_line[0]$_DFFE_PP__155  (.L_HI(net155));
 sg13g2_tiehi \top_inst.sprite_access_inst.sprite_line[10]$_DFFE_PP__156  (.L_HI(net156));
 sg13g2_tiehi \top_inst.sprite_access_inst.sprite_line[11]$_DFFE_PP__157  (.L_HI(net157));
 sg13g2_tiehi \top_inst.sprite_access_inst.sprite_line[1]$_DFFE_PP__158  (.L_HI(net158));
 sg13g2_tiehi \top_inst.sprite_access_inst.sprite_line[2]$_DFFE_PP__159  (.L_HI(net159));
 sg13g2_tiehi \top_inst.sprite_access_inst.sprite_line[3]$_DFFE_PP__160  (.L_HI(net160));
 sg13g2_tiehi \top_inst.sprite_access_inst.sprite_line[4]$_DFFE_PP__161  (.L_HI(net161));
 sg13g2_tiehi \top_inst.sprite_access_inst.sprite_line[5]$_DFFE_PP__162  (.L_HI(net162));
 sg13g2_tiehi \top_inst.sprite_access_inst.sprite_line[6]$_DFFE_PP__163  (.L_HI(net163));
 sg13g2_tiehi \top_inst.sprite_access_inst.sprite_line[7]$_DFFE_PP__164  (.L_HI(net164));
 sg13g2_tiehi \top_inst.sprite_access_inst.sprite_line[8]$_DFFE_PP__165  (.L_HI(net165));
 sg13g2_tiehi \top_inst.sprite_access_inst.sprite_line[9]$_DFFE_PP__166  (.L_HI(net166));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_level_0_1_10_clk (.A(clknet_4_0_0_clk),
    .X(clknet_level_0_1_10_clk));
 sg13g2_buf_2 clkbuf_level_1_1_11_clk (.A(clknet_level_0_1_10_clk),
    .X(clknet_level_1_1_11_clk));
 sg13g2_buf_2 clkbuf_level_2_1_12_clk (.A(clknet_level_1_1_11_clk),
    .X(clknet_level_2_1_12_clk));
 sg13g2_buf_2 clkbuf_level_3_1_13_clk (.A(clknet_level_2_1_12_clk),
    .X(clknet_level_3_1_13_clk));
 sg13g2_buf_2 clkbuf_level_0_1_24_clk (.A(clknet_4_1_0_clk),
    .X(clknet_level_0_1_24_clk));
 sg13g2_buf_2 clkbuf_level_1_1_25_clk (.A(clknet_level_0_1_24_clk),
    .X(clknet_level_1_1_25_clk));
 sg13g2_buf_2 clkbuf_level_2_1_26_clk (.A(clknet_level_1_1_25_clk),
    .X(clknet_level_2_1_26_clk));
 sg13g2_buf_2 clkbuf_level_3_1_27_clk (.A(clknet_level_2_1_26_clk),
    .X(clknet_level_3_1_27_clk));
 sg13g2_buf_2 clkbuf_level_0_1_38_clk (.A(clknet_4_2_0_clk),
    .X(clknet_level_0_1_38_clk));
 sg13g2_buf_2 clkbuf_level_1_1_39_clk (.A(clknet_level_0_1_38_clk),
    .X(clknet_level_1_1_39_clk));
 sg13g2_buf_2 clkbuf_level_2_1_310_clk (.A(clknet_level_1_1_39_clk),
    .X(clknet_level_2_1_310_clk));
 sg13g2_buf_2 clkbuf_level_3_1_311_clk (.A(clknet_level_2_1_310_clk),
    .X(clknet_level_3_1_311_clk));
 sg13g2_buf_2 clkbuf_level_0_1_412_clk (.A(clknet_4_3_0_clk),
    .X(clknet_level_0_1_412_clk));
 sg13g2_buf_2 clkbuf_level_1_1_413_clk (.A(clknet_level_0_1_412_clk),
    .X(clknet_level_1_1_413_clk));
 sg13g2_buf_2 clkbuf_level_2_1_414_clk (.A(clknet_level_1_1_413_clk),
    .X(clknet_level_2_1_414_clk));
 sg13g2_buf_2 clkbuf_level_3_1_415_clk (.A(clknet_level_2_1_414_clk),
    .X(clknet_level_3_1_415_clk));
 sg13g2_buf_2 clkbuf_level_0_1_516_clk (.A(clknet_4_4_0_clk),
    .X(clknet_level_0_1_516_clk));
 sg13g2_buf_2 clkbuf_level_1_1_517_clk (.A(clknet_level_0_1_516_clk),
    .X(clknet_level_1_1_517_clk));
 sg13g2_buf_2 clkbuf_level_2_1_518_clk (.A(clknet_level_1_1_517_clk),
    .X(clknet_level_2_1_518_clk));
 sg13g2_buf_2 clkbuf_level_3_1_519_clk (.A(clknet_level_2_1_518_clk),
    .X(clknet_level_3_1_519_clk));
 sg13g2_buf_2 clkbuf_level_0_1_620_clk (.A(clknet_4_5_0_clk),
    .X(clknet_level_0_1_620_clk));
 sg13g2_buf_2 clkbuf_level_1_1_621_clk (.A(clknet_level_0_1_620_clk),
    .X(clknet_level_1_1_621_clk));
 sg13g2_buf_2 clkbuf_level_2_1_622_clk (.A(clknet_level_1_1_621_clk),
    .X(clknet_level_2_1_622_clk));
 sg13g2_buf_2 clkbuf_level_3_1_623_clk (.A(clknet_level_2_1_622_clk),
    .X(clknet_level_3_1_623_clk));
 sg13g2_buf_2 clkbuf_level_0_1_724_clk (.A(clknet_4_6_0_clk),
    .X(clknet_level_0_1_724_clk));
 sg13g2_buf_2 clkbuf_level_1_1_725_clk (.A(clknet_level_0_1_724_clk),
    .X(clknet_level_1_1_725_clk));
 sg13g2_buf_2 clkbuf_level_2_1_726_clk (.A(clknet_level_1_1_725_clk),
    .X(clknet_level_2_1_726_clk));
 sg13g2_buf_2 clkbuf_level_3_1_727_clk (.A(clknet_level_2_1_726_clk),
    .X(clknet_level_3_1_727_clk));
 sg13g2_buf_2 clkbuf_level_0_1_828_clk (.A(clknet_4_7_0_clk),
    .X(clknet_level_0_1_828_clk));
 sg13g2_buf_2 clkbuf_level_1_1_829_clk (.A(clknet_level_0_1_828_clk),
    .X(clknet_level_1_1_829_clk));
 sg13g2_buf_2 clkbuf_level_2_1_830_clk (.A(clknet_level_1_1_829_clk),
    .X(clknet_level_2_1_830_clk));
 sg13g2_buf_2 clkbuf_level_3_1_831_clk (.A(clknet_level_2_1_830_clk),
    .X(clknet_level_3_1_831_clk));
 sg13g2_buf_2 clkbuf_level_0_1_932_clk (.A(clknet_4_8_0_clk),
    .X(clknet_level_0_1_932_clk));
 sg13g2_buf_2 clkbuf_level_1_1_933_clk (.A(clknet_level_0_1_932_clk),
    .X(clknet_level_1_1_933_clk));
 sg13g2_buf_2 clkbuf_level_2_1_934_clk (.A(clknet_level_1_1_933_clk),
    .X(clknet_level_2_1_934_clk));
 sg13g2_buf_2 clkbuf_level_3_1_935_clk (.A(clknet_level_2_1_934_clk),
    .X(clknet_level_3_1_935_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1036_clk (.A(clknet_4_9_0_clk),
    .X(clknet_level_0_1_1036_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1037_clk (.A(clknet_level_0_1_1036_clk),
    .X(clknet_level_1_1_1037_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1038_clk (.A(clknet_level_1_1_1037_clk),
    .X(clknet_level_2_1_1038_clk));
 sg13g2_buf_2 clkbuf_level_3_1_1039_clk (.A(clknet_level_2_1_1038_clk),
    .X(clknet_level_3_1_1039_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1140_clk (.A(clknet_4_10_0_clk),
    .X(clknet_level_0_1_1140_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1141_clk (.A(clknet_level_0_1_1140_clk),
    .X(clknet_level_1_1_1141_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1142_clk (.A(clknet_level_1_1_1141_clk),
    .X(clknet_level_2_1_1142_clk));
 sg13g2_buf_2 clkbuf_level_3_1_1143_clk (.A(clknet_level_2_1_1142_clk),
    .X(clknet_level_3_1_1143_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1244_clk (.A(clknet_4_11_0_clk),
    .X(clknet_level_0_1_1244_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1245_clk (.A(clknet_level_0_1_1244_clk),
    .X(clknet_level_1_1_1245_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1246_clk (.A(clknet_level_1_1_1245_clk),
    .X(clknet_level_2_1_1246_clk));
 sg13g2_buf_2 clkbuf_level_3_1_1247_clk (.A(clknet_level_2_1_1246_clk),
    .X(clknet_level_3_1_1247_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1348_clk (.A(clknet_4_12_0_clk),
    .X(clknet_level_0_1_1348_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1349_clk (.A(clknet_level_0_1_1348_clk),
    .X(clknet_level_1_1_1349_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1350_clk (.A(clknet_level_1_1_1349_clk),
    .X(clknet_level_2_1_1350_clk));
 sg13g2_buf_2 clkbuf_level_3_1_1351_clk (.A(clknet_level_2_1_1350_clk),
    .X(clknet_level_3_1_1351_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1452_clk (.A(clknet_4_13_0_clk),
    .X(clknet_level_0_1_1452_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1453_clk (.A(clknet_level_0_1_1452_clk),
    .X(clknet_level_1_1_1453_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1454_clk (.A(clknet_level_1_1_1453_clk),
    .X(clknet_level_2_1_1454_clk));
 sg13g2_buf_2 clkbuf_level_3_1_1455_clk (.A(clknet_level_2_1_1454_clk),
    .X(clknet_level_3_1_1455_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1556_clk (.A(clknet_4_14_0_clk),
    .X(clknet_level_0_1_1556_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1557_clk (.A(clknet_level_0_1_1556_clk),
    .X(clknet_level_1_1_1557_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1558_clk (.A(clknet_level_1_1_1557_clk),
    .X(clknet_level_2_1_1558_clk));
 sg13g2_buf_2 clkbuf_level_3_1_1559_clk (.A(clknet_level_2_1_1558_clk),
    .X(clknet_level_3_1_1559_clk));
 sg13g2_buf_2 clkbuf_level_0_1_1660_clk (.A(clknet_4_15_0_clk),
    .X(clknet_level_0_1_1660_clk));
 sg13g2_buf_2 clkbuf_level_1_1_1661_clk (.A(clknet_level_0_1_1660_clk),
    .X(clknet_level_1_1_1661_clk));
 sg13g2_buf_2 clkbuf_level_2_1_1662_clk (.A(clknet_level_1_1_1661_clk),
    .X(clknet_level_2_1_1662_clk));
 sg13g2_buf_2 clkbuf_level_3_1_1663_clk (.A(clknet_level_2_1_1662_clk),
    .X(clknet_level_3_1_1663_clk));
 sg13g2_inv_2 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_inv_2 clkload1 (.A(clknet_4_1_0_clk));
 sg13g2_inv_2 clkload2 (.A(clknet_4_2_0_clk));
 sg13g2_inv_2 clkload3 (.A(clknet_4_3_0_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_4_4_0_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_4_5_0_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_4_6_0_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_4_7_0_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_4_8_0_clk));
 sg13g2_inv_2 clkload9 (.A(clknet_4_9_0_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_4_11_0_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_4_12_0_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_4_13_0_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_4_14_0_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_0__0021_ (.A(_0021_),
    .X(clknet_0__0021_));
 sg13g2_buf_1 clkbuf_1_0__f__0021_ (.A(clknet_0__0021_),
    .X(clknet_1_0__leaf__0021_));
 sg13g2_buf_1 clkbuf_1_1__f__0021_ (.A(clknet_0__0021_),
    .X(clknet_1_1__leaf__0021_));
 sg13g2_buf_1 clkbuf_0__0020_ (.A(_0020_),
    .X(clknet_0__0020_));
 sg13g2_buf_1 clkbuf_1_0__f__0020_ (.A(clknet_0__0020_),
    .X(clknet_1_0__leaf__0020_));
 sg13g2_buf_1 clkbuf_1_1__f__0020_ (.A(clknet_0__0020_),
    .X(clknet_1_1__leaf__0020_));
 sg13g2_buf_1 clkbuf_0__0019_ (.A(_0019_),
    .X(clknet_0__0019_));
 sg13g2_buf_1 clkbuf_1_0__f__0019_ (.A(clknet_0__0019_),
    .X(clknet_1_0__leaf__0019_));
 sg13g2_buf_1 clkbuf_1_1__f__0019_ (.A(clknet_0__0019_),
    .X(clknet_1_1__leaf__0019_));
 sg13g2_buf_1 clkbuf_0__0018_ (.A(_0018_),
    .X(clknet_0__0018_));
 sg13g2_buf_1 clkbuf_1_0__f__0018_ (.A(clknet_0__0018_),
    .X(clknet_1_0__leaf__0018_));
 sg13g2_buf_1 clkbuf_1_1__f__0018_ (.A(clknet_0__0018_),
    .X(clknet_1_1__leaf__0018_));
 sg13g2_buf_1 clkbuf_0__0017_ (.A(_0017_),
    .X(clknet_0__0017_));
 sg13g2_buf_1 clkbuf_1_0__f__0017_ (.A(clknet_0__0017_),
    .X(clknet_1_0__leaf__0017_));
 sg13g2_buf_1 clkbuf_1_1__f__0017_ (.A(clknet_0__0017_),
    .X(clknet_1_1__leaf__0017_));
 sg13g2_buf_1 clkbuf_0__0016_ (.A(_0016_),
    .X(clknet_0__0016_));
 sg13g2_buf_1 clkbuf_1_0__f__0016_ (.A(clknet_0__0016_),
    .X(clknet_1_0__leaf__0016_));
 sg13g2_buf_1 clkbuf_1_1__f__0016_ (.A(clknet_0__0016_),
    .X(clknet_1_1__leaf__0016_));
 sg13g2_buf_1 clkbuf_0__0015_ (.A(_0015_),
    .X(clknet_0__0015_));
 sg13g2_buf_1 clkbuf_1_0__f__0015_ (.A(clknet_0__0015_),
    .X(clknet_1_0__leaf__0015_));
 sg13g2_buf_1 clkbuf_1_1__f__0015_ (.A(clknet_0__0015_),
    .X(clknet_1_1__leaf__0015_));
 sg13g2_buf_1 \clkbuf_0_top_inst.sprite_data_inst.gclk  (.A(\top_inst.sprite_data_inst.gclk ),
    .X(\clknet_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_0_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_0_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_1_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_1_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_2_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_2_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_3_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_3_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_4_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_4_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_5_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_5_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_6_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_6_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_7_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_7_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_8_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_8_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_9_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_9_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_10_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_10_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_11_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_11_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_12_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_12_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_13_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_13_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_14_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_14_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_2 \clkbuf_4_15_0_top_inst.sprite_data_inst.gclk  (.A(\clknet_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_4_15_0_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_0__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_0_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_0__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_1__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_0_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_1__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_2__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_1_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_2__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_3__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_1_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_3__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_4__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_2_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_4__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_5__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_2_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_5__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_6__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_3_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_6__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_7__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_3_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_7__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_8__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_4_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_8__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_9__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_4_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_9__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_10__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_5_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_10__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_11__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_5_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_11__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_12__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_6_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_12__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_13__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_6_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_13__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_14__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_7_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_14__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_15__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_7_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_15__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_16__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_8_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_16__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_17__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_8_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_17__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_18__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_9_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_18__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_19__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_9_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_19__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_20__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_10_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_20__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_21__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_10_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_21__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_22__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_11_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_22__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_23__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_11_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_23__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_24__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_12_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_24__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_25__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_12_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_25__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_26__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_13_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_26__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_27__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_13_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_27__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_28__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_14_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_28__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_29__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_14_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_29__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_30__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_15_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_30__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_buf_1 \clkbuf_5_31__f_top_inst.sprite_data_inst.gclk  (.A(\clknet_4_15_0_top_inst.sprite_data_inst.gclk ),
    .X(\clknet_5_31__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload15 (.A(\clknet_5_1__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload16 (.A(\clknet_5_3__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload17 (.A(\clknet_5_5__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload18 (.A(\clknet_5_7__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload19 (.A(\clknet_5_9__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload20 (.A(\clknet_5_11__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload21 (.A(\clknet_5_13__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload22 (.A(\clknet_5_15__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload23 (.A(\clknet_5_17__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload24 (.A(\clknet_5_19__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload25 (.A(\clknet_5_21__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload26 (.A(\clknet_5_23__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload27 (.A(\clknet_5_25__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload28 (.A(\clknet_5_27__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload29 (.A(\clknet_5_29__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_inv_1 clkload30 (.A(\clknet_5_31__leaf_top_inst.sprite_data_inst.gclk ));
 sg13g2_dlygate4sd3_1 hold1 (.A(\top_inst.spi_mosi_sync ),
    .X(net167));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_fill_2 FILLER_0_35 ();
 sg13g2_fill_1 FILLER_0_37 ();
 sg13g2_fill_1 FILLER_0_64 ();
 sg13g2_fill_1 FILLER_0_68 ();
 sg13g2_fill_1 FILLER_0_95 ();
 sg13g2_fill_1 FILLER_0_99 ();
 sg13g2_decap_4 FILLER_0_152 ();
 sg13g2_fill_1 FILLER_0_156 ();
 sg13g2_fill_1 FILLER_0_313 ();
 sg13g2_decap_4 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_8 FILLER_0_403 ();
 sg13g2_decap_8 FILLER_0_410 ();
 sg13g2_decap_8 FILLER_0_417 ();
 sg13g2_decap_4 FILLER_0_424 ();
 sg13g2_fill_2 FILLER_0_428 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_4 FILLER_1_7 ();
 sg13g2_fill_1 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_44 ();
 sg13g2_decap_4 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_107 ();
 sg13g2_decap_4 FILLER_1_174 ();
 sg13g2_decap_4 FILLER_1_210 ();
 sg13g2_fill_1 FILLER_1_218 ();
 sg13g2_decap_4 FILLER_1_248 ();
 sg13g2_fill_2 FILLER_1_252 ();
 sg13g2_decap_4 FILLER_1_257 ();
 sg13g2_fill_2 FILLER_1_261 ();
 sg13g2_fill_1 FILLER_1_289 ();
 sg13g2_fill_2 FILLER_1_327 ();
 sg13g2_decap_4 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_414 ();
 sg13g2_decap_8 FILLER_1_421 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_decap_4 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_30 ();
 sg13g2_decap_8 FILLER_2_110 ();
 sg13g2_decap_8 FILLER_2_117 ();
 sg13g2_fill_2 FILLER_2_124 ();
 sg13g2_fill_2 FILLER_2_133 ();
 sg13g2_fill_2 FILLER_2_190 ();
 sg13g2_fill_2 FILLER_2_202 ();
 sg13g2_fill_2 FILLER_2_233 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_fill_1 FILLER_2_294 ();
 sg13g2_decap_4 FILLER_2_350 ();
 sg13g2_fill_2 FILLER_2_354 ();
 sg13g2_fill_1 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_416 ();
 sg13g2_decap_8 FILLER_2_423 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_4 FILLER_3_24 ();
 sg13g2_decap_4 FILLER_3_61 ();
 sg13g2_decap_4 FILLER_3_150 ();
 sg13g2_fill_2 FILLER_3_154 ();
 sg13g2_fill_2 FILLER_3_159 ();
 sg13g2_fill_1 FILLER_3_161 ();
 sg13g2_decap_4 FILLER_3_217 ();
 sg13g2_fill_1 FILLER_3_221 ();
 sg13g2_decap_8 FILLER_3_274 ();
 sg13g2_fill_1 FILLER_3_281 ();
 sg13g2_fill_1 FILLER_3_308 ();
 sg13g2_fill_2 FILLER_3_335 ();
 sg13g2_fill_2 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_403 ();
 sg13g2_decap_8 FILLER_3_410 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_4 FILLER_3_424 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_4 FILLER_4_14 ();
 sg13g2_fill_1 FILLER_4_18 ();
 sg13g2_fill_2 FILLER_4_48 ();
 sg13g2_fill_1 FILLER_4_50 ();
 sg13g2_fill_1 FILLER_4_189 ();
 sg13g2_fill_2 FILLER_4_193 ();
 sg13g2_decap_8 FILLER_4_221 ();
 sg13g2_decap_8 FILLER_4_228 ();
 sg13g2_fill_1 FILLER_4_266 ();
 sg13g2_fill_2 FILLER_4_306 ();
 sg13g2_decap_8 FILLER_4_312 ();
 sg13g2_decap_4 FILLER_4_319 ();
 sg13g2_fill_2 FILLER_4_323 ();
 sg13g2_fill_2 FILLER_4_351 ();
 sg13g2_fill_1 FILLER_4_353 ();
 sg13g2_fill_1 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_415 ();
 sg13g2_decap_8 FILLER_4_422 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_39 ();
 sg13g2_fill_1 FILLER_5_46 ();
 sg13g2_decap_8 FILLER_5_73 ();
 sg13g2_decap_8 FILLER_5_80 ();
 sg13g2_fill_1 FILLER_5_100 ();
 sg13g2_decap_8 FILLER_5_160 ();
 sg13g2_fill_2 FILLER_5_171 ();
 sg13g2_fill_2 FILLER_5_202 ();
 sg13g2_fill_2 FILLER_5_238 ();
 sg13g2_fill_1 FILLER_5_240 ();
 sg13g2_fill_2 FILLER_5_282 ();
 sg13g2_fill_1 FILLER_5_284 ();
 sg13g2_decap_8 FILLER_5_311 ();
 sg13g2_decap_8 FILLER_5_318 ();
 sg13g2_decap_4 FILLER_5_328 ();
 sg13g2_decap_4 FILLER_5_370 ();
 sg13g2_fill_2 FILLER_5_374 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_5_409 ();
 sg13g2_decap_8 FILLER_5_416 ();
 sg13g2_decap_8 FILLER_5_423 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_decap_4 FILLER_6_56 ();
 sg13g2_fill_2 FILLER_6_60 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_fill_1 FILLER_6_147 ();
 sg13g2_fill_2 FILLER_6_177 ();
 sg13g2_fill_2 FILLER_6_205 ();
 sg13g2_fill_1 FILLER_6_207 ();
 sg13g2_fill_2 FILLER_6_240 ();
 sg13g2_decap_8 FILLER_6_246 ();
 sg13g2_fill_1 FILLER_6_253 ();
 sg13g2_fill_2 FILLER_6_339 ();
 sg13g2_decap_8 FILLER_6_367 ();
 sg13g2_decap_8 FILLER_6_374 ();
 sg13g2_decap_8 FILLER_6_381 ();
 sg13g2_decap_8 FILLER_6_388 ();
 sg13g2_decap_8 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_6_409 ();
 sg13g2_decap_8 FILLER_6_416 ();
 sg13g2_decap_8 FILLER_6_423 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_4 ();
 sg13g2_fill_1 FILLER_7_31 ();
 sg13g2_fill_2 FILLER_7_35 ();
 sg13g2_fill_1 FILLER_7_37 ();
 sg13g2_fill_2 FILLER_7_72 ();
 sg13g2_fill_1 FILLER_7_74 ();
 sg13g2_fill_1 FILLER_7_104 ();
 sg13g2_fill_1 FILLER_7_131 ();
 sg13g2_fill_1 FILLER_7_184 ();
 sg13g2_fill_2 FILLER_7_216 ();
 sg13g2_fill_1 FILLER_7_218 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_fill_2 FILLER_7_252 ();
 sg13g2_fill_1 FILLER_7_254 ();
 sg13g2_fill_1 FILLER_7_307 ();
 sg13g2_decap_8 FILLER_7_312 ();
 sg13g2_fill_2 FILLER_7_322 ();
 sg13g2_fill_1 FILLER_7_324 ();
 sg13g2_fill_2 FILLER_7_351 ();
 sg13g2_fill_1 FILLER_7_353 ();
 sg13g2_decap_8 FILLER_7_409 ();
 sg13g2_decap_8 FILLER_7_416 ();
 sg13g2_decap_8 FILLER_7_423 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_4 FILLER_8_14 ();
 sg13g2_fill_1 FILLER_8_18 ();
 sg13g2_decap_8 FILLER_8_116 ();
 sg13g2_fill_2 FILLER_8_123 ();
 sg13g2_fill_2 FILLER_8_167 ();
 sg13g2_decap_4 FILLER_8_229 ();
 sg13g2_fill_1 FILLER_8_314 ();
 sg13g2_fill_2 FILLER_8_341 ();
 sg13g2_fill_2 FILLER_8_369 ();
 sg13g2_fill_1 FILLER_8_371 ();
 sg13g2_fill_2 FILLER_8_380 ();
 sg13g2_fill_1 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_decap_4 FILLER_8_424 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_4 FILLER_9_56 ();
 sg13g2_fill_2 FILLER_9_60 ();
 sg13g2_fill_2 FILLER_9_129 ();
 sg13g2_fill_1 FILLER_9_131 ();
 sg13g2_fill_1 FILLER_9_158 ();
 sg13g2_decap_8 FILLER_9_163 ();
 sg13g2_decap_8 FILLER_9_170 ();
 sg13g2_fill_1 FILLER_9_177 ();
 sg13g2_fill_2 FILLER_9_204 ();
 sg13g2_fill_1 FILLER_9_206 ();
 sg13g2_fill_1 FILLER_9_212 ();
 sg13g2_fill_1 FILLER_9_247 ();
 sg13g2_fill_2 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_299 ();
 sg13g2_fill_2 FILLER_9_306 ();
 sg13g2_fill_2 FILLER_9_311 ();
 sg13g2_fill_1 FILLER_9_313 ();
 sg13g2_decap_8 FILLER_9_317 ();
 sg13g2_decap_4 FILLER_9_324 ();
 sg13g2_fill_1 FILLER_9_328 ();
 sg13g2_fill_2 FILLER_9_348 ();
 sg13g2_fill_2 FILLER_9_402 ();
 sg13g2_fill_1 FILLER_9_404 ();
 sg13g2_decap_8 FILLER_9_412 ();
 sg13g2_decap_8 FILLER_9_419 ();
 sg13g2_decap_4 FILLER_9_426 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_fill_1 FILLER_10_70 ();
 sg13g2_fill_1 FILLER_10_79 ();
 sg13g2_fill_1 FILLER_10_87 ();
 sg13g2_fill_2 FILLER_10_114 ();
 sg13g2_fill_1 FILLER_10_171 ();
 sg13g2_fill_2 FILLER_10_198 ();
 sg13g2_fill_1 FILLER_10_200 ();
 sg13g2_fill_1 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_10_409 ();
 sg13g2_decap_8 FILLER_10_416 ();
 sg13g2_decap_8 FILLER_10_423 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_4 FILLER_11_70 ();
 sg13g2_fill_2 FILLER_11_74 ();
 sg13g2_decap_8 FILLER_11_80 ();
 sg13g2_decap_8 FILLER_11_87 ();
 sg13g2_decap_8 FILLER_11_94 ();
 sg13g2_decap_8 FILLER_11_101 ();
 sg13g2_decap_8 FILLER_11_108 ();
 sg13g2_decap_8 FILLER_11_115 ();
 sg13g2_decap_8 FILLER_11_122 ();
 sg13g2_decap_8 FILLER_11_129 ();
 sg13g2_decap_8 FILLER_11_136 ();
 sg13g2_decap_8 FILLER_11_143 ();
 sg13g2_fill_2 FILLER_11_150 ();
 sg13g2_decap_8 FILLER_11_156 ();
 sg13g2_decap_8 FILLER_11_163 ();
 sg13g2_decap_8 FILLER_11_170 ();
 sg13g2_fill_1 FILLER_11_177 ();
 sg13g2_decap_8 FILLER_11_187 ();
 sg13g2_decap_8 FILLER_11_198 ();
 sg13g2_decap_8 FILLER_11_205 ();
 sg13g2_decap_8 FILLER_11_212 ();
 sg13g2_decap_8 FILLER_11_219 ();
 sg13g2_decap_8 FILLER_11_226 ();
 sg13g2_decap_8 FILLER_11_233 ();
 sg13g2_decap_8 FILLER_11_240 ();
 sg13g2_fill_2 FILLER_11_247 ();
 sg13g2_fill_1 FILLER_11_249 ();
 sg13g2_fill_2 FILLER_11_254 ();
 sg13g2_fill_2 FILLER_11_259 ();
 sg13g2_fill_1 FILLER_11_261 ();
 sg13g2_decap_4 FILLER_11_293 ();
 sg13g2_fill_2 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_403 ();
 sg13g2_decap_8 FILLER_11_410 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_4 FILLER_11_424 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_4 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_166 ();
 sg13g2_fill_1 FILLER_12_173 ();
 sg13g2_fill_1 FILLER_12_196 ();
 sg13g2_fill_1 FILLER_12_202 ();
 sg13g2_fill_1 FILLER_12_226 ();
 sg13g2_fill_1 FILLER_12_253 ();
 sg13g2_decap_4 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_292 ();
 sg13g2_fill_2 FILLER_12_299 ();
 sg13g2_decap_8 FILLER_12_311 ();
 sg13g2_decap_4 FILLER_12_318 ();
 sg13g2_fill_2 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_353 ();
 sg13g2_fill_2 FILLER_12_360 ();
 sg13g2_fill_1 FILLER_12_362 ();
 sg13g2_decap_8 FILLER_12_373 ();
 sg13g2_decap_8 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_4 FILLER_12_394 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_fill_2 FILLER_13_105 ();
 sg13g2_fill_1 FILLER_13_107 ();
 sg13g2_decap_4 FILLER_13_139 ();
 sg13g2_fill_1 FILLER_13_143 ();
 sg13g2_fill_1 FILLER_13_202 ();
 sg13g2_fill_1 FILLER_13_208 ();
 sg13g2_decap_8 FILLER_13_226 ();
 sg13g2_fill_2 FILLER_13_233 ();
 sg13g2_fill_1 FILLER_13_254 ();
 sg13g2_fill_1 FILLER_13_267 ();
 sg13g2_fill_1 FILLER_13_273 ();
 sg13g2_fill_1 FILLER_13_279 ();
 sg13g2_fill_2 FILLER_13_311 ();
 sg13g2_fill_1 FILLER_13_313 ();
 sg13g2_decap_4 FILLER_13_340 ();
 sg13g2_fill_1 FILLER_13_344 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_4 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_411 ();
 sg13g2_decap_8 FILLER_13_418 ();
 sg13g2_decap_4 FILLER_13_425 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_4 FILLER_14_105 ();
 sg13g2_fill_1 FILLER_14_109 ();
 sg13g2_decap_4 FILLER_14_115 ();
 sg13g2_fill_1 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_134 ();
 sg13g2_decap_8 FILLER_14_141 ();
 sg13g2_fill_1 FILLER_14_148 ();
 sg13g2_fill_2 FILLER_14_152 ();
 sg13g2_fill_1 FILLER_14_154 ();
 sg13g2_fill_2 FILLER_14_159 ();
 sg13g2_fill_2 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_230 ();
 sg13g2_fill_1 FILLER_14_237 ();
 sg13g2_fill_1 FILLER_14_255 ();
 sg13g2_fill_2 FILLER_14_293 ();
 sg13g2_decap_4 FILLER_14_309 ();
 sg13g2_fill_1 FILLER_14_313 ();
 sg13g2_fill_2 FILLER_14_366 ();
 sg13g2_fill_1 FILLER_14_398 ();
 sg13g2_decap_8 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_14_412 ();
 sg13g2_decap_8 FILLER_14_419 ();
 sg13g2_decap_4 FILLER_14_426 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_fill_2 FILLER_15_91 ();
 sg13g2_decap_4 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_159 ();
 sg13g2_fill_1 FILLER_15_173 ();
 sg13g2_fill_1 FILLER_15_178 ();
 sg13g2_fill_1 FILLER_15_186 ();
 sg13g2_fill_2 FILLER_15_192 ();
 sg13g2_decap_4 FILLER_15_199 ();
 sg13g2_fill_1 FILLER_15_203 ();
 sg13g2_fill_2 FILLER_15_235 ();
 sg13g2_decap_4 FILLER_15_241 ();
 sg13g2_fill_1 FILLER_15_300 ();
 sg13g2_decap_4 FILLER_15_327 ();
 sg13g2_fill_1 FILLER_15_331 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_fill_2 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_4 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_22 ();
 sg13g2_decap_4 FILLER_16_29 ();
 sg13g2_decap_8 FILLER_16_40 ();
 sg13g2_fill_2 FILLER_16_47 ();
 sg13g2_fill_2 FILLER_16_53 ();
 sg13g2_fill_1 FILLER_16_55 ();
 sg13g2_decap_8 FILLER_16_95 ();
 sg13g2_fill_2 FILLER_16_102 ();
 sg13g2_decap_4 FILLER_16_116 ();
 sg13g2_fill_2 FILLER_16_130 ();
 sg13g2_fill_1 FILLER_16_158 ();
 sg13g2_fill_1 FILLER_16_200 ();
 sg13g2_fill_1 FILLER_16_235 ();
 sg13g2_fill_2 FILLER_16_241 ();
 sg13g2_fill_1 FILLER_16_243 ();
 sg13g2_fill_1 FILLER_16_260 ();
 sg13g2_fill_2 FILLER_16_266 ();
 sg13g2_fill_1 FILLER_16_268 ();
 sg13g2_fill_2 FILLER_16_274 ();
 sg13g2_fill_2 FILLER_16_323 ();
 sg13g2_fill_1 FILLER_16_338 ();
 sg13g2_fill_1 FILLER_16_344 ();
 sg13g2_fill_1 FILLER_16_353 ();
 sg13g2_fill_2 FILLER_16_362 ();
 sg13g2_fill_1 FILLER_16_364 ();
 sg13g2_fill_2 FILLER_16_370 ();
 sg13g2_fill_1 FILLER_16_372 ();
 sg13g2_decap_8 FILLER_16_409 ();
 sg13g2_decap_8 FILLER_16_416 ();
 sg13g2_decap_8 FILLER_16_423 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_fill_2 FILLER_17_11 ();
 sg13g2_fill_2 FILLER_17_69 ();
 sg13g2_fill_2 FILLER_17_117 ();
 sg13g2_fill_1 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_160 ();
 sg13g2_fill_2 FILLER_17_166 ();
 sg13g2_fill_2 FILLER_17_173 ();
 sg13g2_fill_2 FILLER_17_179 ();
 sg13g2_fill_2 FILLER_17_186 ();
 sg13g2_fill_2 FILLER_17_219 ();
 sg13g2_fill_2 FILLER_17_238 ();
 sg13g2_fill_1 FILLER_17_240 ();
 sg13g2_fill_2 FILLER_17_344 ();
 sg13g2_fill_1 FILLER_17_350 ();
 sg13g2_fill_2 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_17_412 ();
 sg13g2_decap_8 FILLER_17_419 ();
 sg13g2_decap_4 FILLER_17_426 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_36 ();
 sg13g2_fill_1 FILLER_18_59 ();
 sg13g2_fill_1 FILLER_18_65 ();
 sg13g2_fill_2 FILLER_18_71 ();
 sg13g2_fill_1 FILLER_18_73 ();
 sg13g2_fill_2 FILLER_18_82 ();
 sg13g2_fill_2 FILLER_18_89 ();
 sg13g2_fill_1 FILLER_18_91 ();
 sg13g2_fill_2 FILLER_18_142 ();
 sg13g2_fill_1 FILLER_18_197 ();
 sg13g2_fill_1 FILLER_18_234 ();
 sg13g2_fill_2 FILLER_18_239 ();
 sg13g2_fill_2 FILLER_18_245 ();
 sg13g2_fill_1 FILLER_18_283 ();
 sg13g2_fill_1 FILLER_18_306 ();
 sg13g2_fill_1 FILLER_18_311 ();
 sg13g2_fill_1 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_417 ();
 sg13g2_decap_4 FILLER_18_424 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_fill_2 FILLER_19_39 ();
 sg13g2_fill_2 FILLER_19_48 ();
 sg13g2_fill_1 FILLER_19_50 ();
 sg13g2_fill_2 FILLER_19_130 ();
 sg13g2_fill_1 FILLER_19_132 ();
 sg13g2_fill_2 FILLER_19_160 ();
 sg13g2_fill_1 FILLER_19_173 ();
 sg13g2_decap_8 FILLER_19_194 ();
 sg13g2_decap_4 FILLER_19_201 ();
 sg13g2_fill_2 FILLER_19_222 ();
 sg13g2_fill_1 FILLER_19_233 ();
 sg13g2_fill_2 FILLER_19_264 ();
 sg13g2_fill_2 FILLER_19_292 ();
 sg13g2_fill_1 FILLER_19_299 ();
 sg13g2_decap_8 FILLER_19_383 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_fill_1 FILLER_20_56 ();
 sg13g2_fill_2 FILLER_20_84 ();
 sg13g2_fill_2 FILLER_20_98 ();
 sg13g2_fill_1 FILLER_20_100 ();
 sg13g2_fill_2 FILLER_20_131 ();
 sg13g2_fill_1 FILLER_20_133 ();
 sg13g2_fill_2 FILLER_20_160 ();
 sg13g2_fill_1 FILLER_20_170 ();
 sg13g2_fill_2 FILLER_20_183 ();
 sg13g2_fill_1 FILLER_20_185 ();
 sg13g2_fill_2 FILLER_20_195 ();
 sg13g2_fill_2 FILLER_20_228 ();
 sg13g2_fill_2 FILLER_20_277 ();
 sg13g2_fill_2 FILLER_20_283 ();
 sg13g2_fill_2 FILLER_20_316 ();
 sg13g2_fill_2 FILLER_20_328 ();
 sg13g2_fill_1 FILLER_20_330 ();
 sg13g2_fill_1 FILLER_20_346 ();
 sg13g2_fill_1 FILLER_20_370 ();
 sg13g2_fill_1 FILLER_20_401 ();
 sg13g2_decap_8 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_20_414 ();
 sg13g2_decap_8 FILLER_20_421 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_fill_2 FILLER_21_61 ();
 sg13g2_fill_2 FILLER_21_84 ();
 sg13g2_fill_1 FILLER_21_86 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_fill_2 FILLER_21_100 ();
 sg13g2_fill_1 FILLER_21_102 ();
 sg13g2_fill_2 FILLER_21_133 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_fill_1 FILLER_21_169 ();
 sg13g2_fill_1 FILLER_21_187 ();
 sg13g2_fill_1 FILLER_21_194 ();
 sg13g2_fill_2 FILLER_21_203 ();
 sg13g2_fill_2 FILLER_21_209 ();
 sg13g2_fill_2 FILLER_21_215 ();
 sg13g2_fill_2 FILLER_21_221 ();
 sg13g2_decap_4 FILLER_21_228 ();
 sg13g2_decap_4 FILLER_21_237 ();
 sg13g2_decap_4 FILLER_21_268 ();
 sg13g2_fill_2 FILLER_21_272 ();
 sg13g2_fill_1 FILLER_21_286 ();
 sg13g2_fill_1 FILLER_21_292 ();
 sg13g2_fill_1 FILLER_21_298 ();
 sg13g2_fill_2 FILLER_21_303 ();
 sg13g2_decap_4 FILLER_21_313 ();
 sg13g2_fill_1 FILLER_21_317 ();
 sg13g2_fill_1 FILLER_21_322 ();
 sg13g2_fill_1 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_422 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_22 ();
 sg13g2_fill_1 FILLER_22_96 ();
 sg13g2_fill_1 FILLER_22_111 ();
 sg13g2_fill_1 FILLER_22_117 ();
 sg13g2_fill_2 FILLER_22_158 ();
 sg13g2_fill_2 FILLER_22_163 ();
 sg13g2_fill_1 FILLER_22_248 ();
 sg13g2_fill_2 FILLER_22_280 ();
 sg13g2_fill_2 FILLER_22_291 ();
 sg13g2_fill_1 FILLER_22_340 ();
 sg13g2_fill_2 FILLER_22_345 ();
 sg13g2_fill_2 FILLER_22_360 ();
 sg13g2_decap_4 FILLER_22_398 ();
 sg13g2_fill_1 FILLER_22_402 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_fill_2 FILLER_23_34 ();
 sg13g2_fill_1 FILLER_23_36 ();
 sg13g2_fill_1 FILLER_23_94 ();
 sg13g2_fill_1 FILLER_23_104 ();
 sg13g2_fill_1 FILLER_23_115 ();
 sg13g2_fill_2 FILLER_23_131 ();
 sg13g2_fill_1 FILLER_23_138 ();
 sg13g2_decap_4 FILLER_23_152 ();
 sg13g2_fill_1 FILLER_23_163 ();
 sg13g2_decap_4 FILLER_23_199 ();
 sg13g2_fill_1 FILLER_23_203 ();
 sg13g2_fill_1 FILLER_23_208 ();
 sg13g2_fill_1 FILLER_23_213 ();
 sg13g2_fill_1 FILLER_23_219 ();
 sg13g2_fill_1 FILLER_23_267 ();
 sg13g2_fill_1 FILLER_23_281 ();
 sg13g2_fill_2 FILLER_23_316 ();
 sg13g2_decap_8 FILLER_23_421 ();
 sg13g2_fill_2 FILLER_23_428 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_15 ();
 sg13g2_fill_1 FILLER_24_26 ();
 sg13g2_fill_1 FILLER_24_61 ();
 sg13g2_fill_1 FILLER_24_97 ();
 sg13g2_fill_2 FILLER_24_183 ();
 sg13g2_fill_1 FILLER_24_192 ();
 sg13g2_fill_2 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_205 ();
 sg13g2_fill_2 FILLER_24_219 ();
 sg13g2_fill_2 FILLER_24_250 ();
 sg13g2_fill_1 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_268 ();
 sg13g2_fill_2 FILLER_24_275 ();
 sg13g2_fill_1 FILLER_24_372 ();
 sg13g2_fill_1 FILLER_24_399 ();
 sg13g2_fill_1 FILLER_25_51 ();
 sg13g2_fill_1 FILLER_25_67 ();
 sg13g2_fill_2 FILLER_25_73 ();
 sg13g2_fill_2 FILLER_25_114 ();
 sg13g2_fill_2 FILLER_25_205 ();
 sg13g2_fill_1 FILLER_25_207 ();
 sg13g2_decap_8 FILLER_25_221 ();
 sg13g2_fill_1 FILLER_25_239 ();
 sg13g2_fill_2 FILLER_25_283 ();
 sg13g2_fill_1 FILLER_25_285 ();
 sg13g2_decap_8 FILLER_25_296 ();
 sg13g2_fill_2 FILLER_25_303 ();
 sg13g2_fill_1 FILLER_25_310 ();
 sg13g2_fill_1 FILLER_25_320 ();
 sg13g2_fill_1 FILLER_25_326 ();
 sg13g2_fill_1 FILLER_25_337 ();
 sg13g2_fill_2 FILLER_25_343 ();
 sg13g2_fill_2 FILLER_25_376 ();
 sg13g2_fill_1 FILLER_25_403 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_fill_2 FILLER_25_427 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_51 ();
 sg13g2_fill_1 FILLER_26_87 ();
 sg13g2_decap_4 FILLER_26_183 ();
 sg13g2_fill_2 FILLER_26_204 ();
 sg13g2_decap_8 FILLER_26_220 ();
 sg13g2_fill_2 FILLER_26_227 ();
 sg13g2_fill_1 FILLER_26_229 ();
 sg13g2_fill_2 FILLER_26_240 ();
 sg13g2_fill_1 FILLER_26_250 ();
 sg13g2_decap_8 FILLER_26_268 ();
 sg13g2_fill_1 FILLER_26_275 ();
 sg13g2_fill_1 FILLER_26_280 ();
 sg13g2_fill_1 FILLER_26_289 ();
 sg13g2_fill_1 FILLER_26_298 ();
 sg13g2_fill_1 FILLER_26_304 ();
 sg13g2_fill_1 FILLER_26_310 ();
 sg13g2_fill_2 FILLER_26_316 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_fill_1 FILLER_26_388 ();
 sg13g2_fill_2 FILLER_26_411 ();
 sg13g2_fill_1 FILLER_26_413 ();
 sg13g2_fill_2 FILLER_26_418 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_20 ();
 sg13g2_fill_1 FILLER_27_22 ();
 sg13g2_fill_2 FILLER_27_38 ();
 sg13g2_fill_2 FILLER_27_60 ();
 sg13g2_fill_1 FILLER_27_100 ();
 sg13g2_fill_1 FILLER_27_111 ();
 sg13g2_fill_1 FILLER_27_117 ();
 sg13g2_fill_1 FILLER_27_134 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_165 ();
 sg13g2_fill_1 FILLER_27_181 ();
 sg13g2_decap_8 FILLER_27_225 ();
 sg13g2_fill_1 FILLER_27_256 ();
 sg13g2_decap_8 FILLER_27_264 ();
 sg13g2_fill_1 FILLER_27_326 ();
 sg13g2_fill_1 FILLER_27_331 ();
 sg13g2_fill_2 FILLER_27_394 ();
 sg13g2_fill_1 FILLER_28_47 ();
 sg13g2_fill_1 FILLER_28_97 ();
 sg13g2_fill_2 FILLER_28_130 ();
 sg13g2_fill_1 FILLER_28_132 ();
 sg13g2_fill_1 FILLER_28_157 ();
 sg13g2_fill_2 FILLER_28_163 ();
 sg13g2_decap_8 FILLER_28_256 ();
 sg13g2_fill_2 FILLER_28_276 ();
 sg13g2_fill_1 FILLER_28_278 ();
 sg13g2_fill_1 FILLER_28_305 ();
 sg13g2_fill_1 FILLER_28_322 ();
 sg13g2_decap_4 FILLER_28_327 ();
 sg13g2_fill_2 FILLER_28_376 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_23 ();
 sg13g2_fill_1 FILLER_29_94 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_121 ();
 sg13g2_fill_1 FILLER_29_142 ();
 sg13g2_fill_1 FILLER_29_167 ();
 sg13g2_fill_1 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_203 ();
 sg13g2_decap_4 FILLER_29_247 ();
 sg13g2_fill_2 FILLER_29_258 ();
 sg13g2_fill_2 FILLER_29_284 ();
 sg13g2_fill_2 FILLER_29_315 ();
 sg13g2_fill_1 FILLER_29_317 ();
 sg13g2_fill_1 FILLER_29_329 ();
 sg13g2_fill_1 FILLER_29_335 ();
 sg13g2_fill_2 FILLER_29_342 ();
 sg13g2_fill_2 FILLER_29_350 ();
 sg13g2_fill_1 FILLER_29_356 ();
 sg13g2_fill_1 FILLER_29_363 ();
 sg13g2_fill_1 FILLER_29_369 ();
 sg13g2_fill_1 FILLER_29_380 ();
 sg13g2_fill_2 FILLER_29_415 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_28 ();
 sg13g2_fill_2 FILLER_30_60 ();
 sg13g2_fill_1 FILLER_30_62 ();
 sg13g2_fill_2 FILLER_30_100 ();
 sg13g2_fill_1 FILLER_30_146 ();
 sg13g2_fill_2 FILLER_30_219 ();
 sg13g2_fill_2 FILLER_30_240 ();
 sg13g2_fill_2 FILLER_30_247 ();
 sg13g2_fill_2 FILLER_30_304 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_fill_1 FILLER_30_325 ();
 sg13g2_fill_2 FILLER_30_343 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_56 ();
 sg13g2_fill_2 FILLER_31_67 ();
 sg13g2_fill_1 FILLER_31_90 ();
 sg13g2_fill_2 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_fill_1 FILLER_31_173 ();
 sg13g2_fill_2 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_241 ();
 sg13g2_fill_1 FILLER_31_282 ();
 sg13g2_fill_2 FILLER_31_294 ();
 sg13g2_fill_1 FILLER_31_296 ();
 sg13g2_fill_2 FILLER_31_302 ();
 sg13g2_fill_1 FILLER_31_304 ();
 sg13g2_fill_2 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_350 ();
 sg13g2_fill_1 FILLER_32_34 ();
 sg13g2_fill_2 FILLER_32_55 ();
 sg13g2_fill_1 FILLER_32_57 ();
 sg13g2_fill_2 FILLER_32_170 ();
 sg13g2_fill_1 FILLER_32_172 ();
 sg13g2_fill_2 FILLER_32_193 ();
 sg13g2_fill_2 FILLER_32_199 ();
 sg13g2_fill_2 FILLER_32_241 ();
 sg13g2_fill_1 FILLER_32_265 ();
 sg13g2_fill_2 FILLER_32_302 ();
 sg13g2_fill_2 FILLER_32_356 ();
 sg13g2_fill_2 FILLER_32_363 ();
 sg13g2_fill_2 FILLER_32_391 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_82 ();
 sg13g2_fill_1 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_115 ();
 sg13g2_fill_1 FILLER_33_166 ();
 sg13g2_fill_1 FILLER_33_191 ();
 sg13g2_fill_1 FILLER_33_217 ();
 sg13g2_fill_2 FILLER_33_246 ();
 sg13g2_fill_1 FILLER_33_266 ();
 sg13g2_fill_1 FILLER_33_274 ();
 sg13g2_fill_1 FILLER_33_291 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_fill_1 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_371 ();
 sg13g2_fill_1 FILLER_33_387 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_27 ();
 sg13g2_fill_2 FILLER_34_140 ();
 sg13g2_fill_2 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_149 ();
 sg13g2_fill_1 FILLER_34_166 ();
 sg13g2_fill_1 FILLER_34_183 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_2 FILLER_34_205 ();
 sg13g2_fill_2 FILLER_34_254 ();
 sg13g2_fill_2 FILLER_34_296 ();
 sg13g2_fill_2 FILLER_34_345 ();
 sg13g2_fill_2 FILLER_34_380 ();
 sg13g2_fill_1 FILLER_34_402 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_fill_1 FILLER_35_44 ();
 sg13g2_fill_2 FILLER_35_50 ();
 sg13g2_fill_1 FILLER_35_105 ();
 sg13g2_fill_1 FILLER_35_121 ();
 sg13g2_fill_1 FILLER_35_137 ();
 sg13g2_fill_2 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_149 ();
 sg13g2_fill_2 FILLER_35_166 ();
 sg13g2_fill_1 FILLER_35_188 ();
 sg13g2_fill_1 FILLER_35_194 ();
 sg13g2_fill_2 FILLER_35_313 ();
 sg13g2_fill_1 FILLER_35_324 ();
 sg13g2_fill_2 FILLER_35_355 ();
 sg13g2_fill_2 FILLER_35_422 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_9 ();
 sg13g2_fill_2 FILLER_36_122 ();
 sg13g2_fill_1 FILLER_36_124 ();
 sg13g2_fill_1 FILLER_36_144 ();
 sg13g2_fill_2 FILLER_36_161 ();
 sg13g2_fill_1 FILLER_36_163 ();
 sg13g2_fill_1 FILLER_36_270 ();
 sg13g2_fill_2 FILLER_36_276 ();
 sg13g2_fill_2 FILLER_36_283 ();
 sg13g2_fill_2 FILLER_36_289 ();
 sg13g2_fill_2 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_355 ();
 sg13g2_fill_2 FILLER_36_392 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_fill_2 FILLER_37_109 ();
 sg13g2_fill_1 FILLER_37_111 ();
 sg13g2_fill_2 FILLER_37_127 ();
 sg13g2_fill_2 FILLER_37_134 ();
 sg13g2_fill_1 FILLER_37_136 ();
 sg13g2_fill_2 FILLER_37_153 ();
 sg13g2_fill_1 FILLER_37_275 ();
 sg13g2_fill_2 FILLER_37_284 ();
 sg13g2_fill_2 FILLER_37_360 ();
 sg13g2_fill_2 FILLER_37_402 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_54 ();
 sg13g2_fill_2 FILLER_38_73 ();
 sg13g2_fill_2 FILLER_38_80 ();
 sg13g2_fill_1 FILLER_38_82 ();
 sg13g2_fill_2 FILLER_38_129 ();
 sg13g2_fill_1 FILLER_38_131 ();
 sg13g2_fill_1 FILLER_38_141 ();
 sg13g2_fill_1 FILLER_38_277 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_fill_1 FILLER_38_327 ();
endmodule
